--------------------------------------------------------------------------------
--                         ModuloCounter_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_13_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 12 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid310732
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid310732 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid310732 is
signal XX_m310733 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m310733 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m310733 <= X ;
   YY_m310733 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid310736
--                   (IntAdderClassical_33_f500_uid310738)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid310736 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid310736 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid310732 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid310736 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid310732  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid310736  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_13_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid311803_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid311805)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid311803_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid311803_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid311808
--                  (IntAdderAlternative_27_f250_uid311812)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid311808 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid311808 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid311815
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid311815 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid311815 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid311818
--                   (IntAdderClassical_34_f250_uid311820)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid311818 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid311818 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid311803
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid311803 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid311803 is
   component FPAdd_8_23_uid311803_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid311808 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid311815 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid311818 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid311803_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid311808  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid311815  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid311818  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid311803 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid311803  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_8_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
         iS_7 when "111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_11_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_11_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_11_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_12_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid312606_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid312608)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid312606_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid312606_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid312611
--                  (IntAdderAlternative_27_f250_uid312615)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid312611 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid312611 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid312618
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid312618 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid312618 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid312621
--                   (IntAdderClassical_34_f250_uid312623)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid312621 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid312621 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid312606
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid312606 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid312606 is
   component FPAdd_8_23_uid312606_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid312611 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid312618 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid312621 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid312606_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid312611  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid312618  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid312621  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid312606 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid312606  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_4_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
         iS_3 when "11",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_7_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 81 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      Y <= s80;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 54 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      Y <= s53;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 52 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      Y <= s51;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      Y <= s62;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 50 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      Y <= s49;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 48 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      Y <= s47;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 76 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      Y <= s75;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 42 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      Y <= s41;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 66 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      Y <= s65;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 51 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      Y <= s50;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "000" when "0111",
      "110" when "1000",
      "010" when "1001",
      "001" when "1010",
      "111" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "111" when "0111",
      "100" when "1000",
      "010" when "1001",
      "001" when "1010",
      "110" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0001" when "0000",
      "0110" when "0001",
      "1010" when "0010",
      "1001" when "0011",
      "0000" when "0100",
      "0000" when "0101",
      "0000" when "0110",
      "0101" when "0111",
      "0011" when "1000",
      "1000" when "1001",
      "0111" when "1010",
      "0010" when "1011",
      "0100" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0001" when "0000",
      "0000" when "0001",
      "1000" when "0010",
      "0111" when "0011",
      "0000" when "0100",
      "1010" when "0101",
      "0000" when "0110",
      "1001" when "0111",
      "0010" when "1000",
      "0110" when "1001",
      "0100" when "1010",
      "0101" when "1011",
      "0011" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0110" when "0001",
      "0100" when "0010",
      "0101" when "0011",
      "0000" when "0100",
      "0010" when "0101",
      "1000" when "0110",
      "1010" when "0111",
      "0111" when "1000",
      "0011" when "1001",
      "1001" when "1010",
      "1011" when "1011",
      "0001" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0110" when "0001",
      "1010" when "0010",
      "1011" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1001" when "0110",
      "0011" when "0111",
      "0111" when "1000",
      "0010" when "1001",
      "1000" when "1010",
      "0100" when "1011",
      "0101" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "010" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "101" when "0101",
      "000" when "0110",
      "000" when "0111",
      "111" when "1000",
      "011" when "1001",
      "100" when "1010",
      "001" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "010" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "111" when "0111",
      "000" when "1000",
      "101" when "1001",
      "100" when "1010",
      "001" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "00" when "0001",
      "00" when "0010",
      "10" when "0011",
      "00" when "0100",
      "11" when "0101",
      "01" when "0110",
      "00" when "0111",
      "00" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when "1100",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "00" when "0001",
      "00" when "0010",
      "10" when "0011",
      "00" when "0100",
      "11" when "0101",
      "01" when "0110",
      "00" when "0111",
      "00" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when "1100",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "100" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "010" when "0000",
      "001" when "0001",
      "000" when "0010",
      "110" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "100" when "0111",
      "000" when "1000",
      "101" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 86 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      Y <= s85;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 69 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      Y <= s68;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 55 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      Y <= s54;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 62 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      Y <= s61;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 59 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      Y <= s58;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 40 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      Y <= s39;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 67 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      Y <= s66;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      Y <= s40;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 64 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      Y <= s63;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 45 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      Y <= s44;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      Y <= s32;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 99 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      Y <= s98;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_3 : in std_logic_vector(31 downto 0);
          R_U_0 : in std_logic_vector(31 downto 0);
          R_U_1 : in std_logic_vector(31 downto 0);
          R_U_2 : in std_logic_vector(31 downto 0);
          R_U_3 : in std_logic_vector(31 downto 0);
          R_V_0 : in std_logic_vector(31 downto 0);
          R_V_1 : in std_logic_vector(31 downto 0);
          R_V_2 : in std_logic_vector(31 downto 0);
          R_V_3 : in std_logic_vector(31 downto 0);
          R_W_0 : in std_logic_vector(31 downto 0);
          R_W_1 : in std_logic_vector(31 downto 0);
          R_W_2 : in std_logic_vector(31 downto 0);
          R_W_3 : in std_logic_vector(31 downto 0);
          Inv_11_0 : out std_logic_vector(31 downto 0);
          Inv_11_1 : out std_logic_vector(31 downto 0);
          Inv_11_2 : out std_logic_vector(31 downto 0);
          Inv_11_3 : out std_logic_vector(31 downto 0);
          Inv_12_0 : out std_logic_vector(31 downto 0);
          Inv_12_1 : out std_logic_vector(31 downto 0);
          Inv_12_2 : out std_logic_vector(31 downto 0);
          Inv_12_3 : out std_logic_vector(31 downto 0);
          Inv_13_0 : out std_logic_vector(31 downto 0);
          Inv_13_1 : out std_logic_vector(31 downto 0);
          Inv_13_2 : out std_logic_vector(31 downto 0);
          Inv_13_3 : out std_logic_vector(31 downto 0);
          Inv_21_0 : out std_logic_vector(31 downto 0);
          Inv_21_1 : out std_logic_vector(31 downto 0);
          Inv_21_2 : out std_logic_vector(31 downto 0);
          Inv_21_3 : out std_logic_vector(31 downto 0);
          Inv_22_0 : out std_logic_vector(31 downto 0);
          Inv_22_1 : out std_logic_vector(31 downto 0);
          Inv_22_2 : out std_logic_vector(31 downto 0);
          Inv_22_3 : out std_logic_vector(31 downto 0);
          Inv_23_0 : out std_logic_vector(31 downto 0);
          Inv_23_1 : out std_logic_vector(31 downto 0);
          Inv_23_2 : out std_logic_vector(31 downto 0);
          Inv_23_3 : out std_logic_vector(31 downto 0);
          Inv_31_0 : out std_logic_vector(31 downto 0);
          Inv_31_1 : out std_logic_vector(31 downto 0);
          Inv_31_2 : out std_logic_vector(31 downto 0);
          Inv_31_3 : out std_logic_vector(31 downto 0);
          Inv_32_0 : out std_logic_vector(31 downto 0);
          Inv_32_1 : out std_logic_vector(31 downto 0);
          Inv_32_2 : out std_logic_vector(31 downto 0);
          Inv_32_3 : out std_logic_vector(31 downto 0);
          Inv_33_0 : out std_logic_vector(31 downto 0);
          Inv_33_1 : out std_logic_vector(31 downto 0);
          Inv_33_2 : out std_logic_vector(31 downto 0);
          Inv_33_3 : out std_logic_vector(31 downto 0);
          Inv_41_0 : out std_logic_vector(31 downto 0);
          Inv_41_1 : out std_logic_vector(31 downto 0);
          Inv_41_2 : out std_logic_vector(31 downto 0);
          Inv_41_3 : out std_logic_vector(31 downto 0);
          Inv_42_0 : out std_logic_vector(31 downto 0);
          Inv_42_1 : out std_logic_vector(31 downto 0);
          Inv_42_2 : out std_logic_vector(31 downto 0);
          Inv_42_3 : out std_logic_vector(31 downto 0);
          Inv_43_0 : out std_logic_vector(31 downto 0);
          Inv_43_1 : out std_logic_vector(31 downto 0);
          Inv_43_2 : out std_logic_vector(31 downto 0);
          Inv_43_3 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_13_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_13_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_8_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_11_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_12_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_4_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_7_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount131_out : std_logic_vector(3 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add17_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add17_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add17_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product103_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product103_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product103_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product103_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product103_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product103_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product106_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product106_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product106_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product107_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product107_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product107_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product181_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product461_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product911_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product97_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product97_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product97_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract1_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay40No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay58No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay99No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay101No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay56No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay50No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay86No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_3_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add121_3_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add22_3_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add22_3_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product97_3_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product97_3_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add10_3_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add10_3_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product3_3_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product3_3_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No6_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No7_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No2_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No4_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No4_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No6_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No3_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No2_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No6_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay58No1_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No8_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No4_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay101No_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No1_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No5_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No4_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay99No1_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No2_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No7_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay86No6_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No6_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No4_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No9_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No1_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No6_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No3_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No2_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No7_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No15_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No2_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No128_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No1_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay56No3_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No41_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No3_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No1_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No2_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No2_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No8_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay85No5_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No7_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No2_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No8_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No10_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No4_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No5_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No7_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Add141_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Add141_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Add17_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Add17_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay98No1_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Add22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Add22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No9_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No3_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No5_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay108No2_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product113_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product113_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No4_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay54No_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No1_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product103_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product103_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No5_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No1_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product103_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product103_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No7_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No6_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No3_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product106_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product106_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No1_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product107_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product107_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No9_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product181_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product181_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product461_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product461_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product68_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product68_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product911_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product911_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product97_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product97_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No10_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay50No_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No1_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay40No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Add10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Add10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No16_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No1_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount131_instance: ModuloCounter_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount131_out);
Ldiff_UU_del_1_0_IEEE <= Ldiff_UU_del_1_0;
   Ldiff_UU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_0_out,
                 X => Ldiff_UU_del_1_0_IEEE);
Ldiff_UU_del_1_1_IEEE <= Ldiff_UU_del_1_1;
   Ldiff_UU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_1_out,
                 X => Ldiff_UU_del_1_1_IEEE);
Ldiff_UU_del_1_2_IEEE <= Ldiff_UU_del_1_2;
   Ldiff_UU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_2_out,
                 X => Ldiff_UU_del_1_2_IEEE);
Ldiff_UU_del_1_3_IEEE <= Ldiff_UU_del_1_3;
   Ldiff_UU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_3_out,
                 X => Ldiff_UU_del_1_3_IEEE);
Ldiff_UV_del_1_0_IEEE <= Ldiff_UV_del_1_0;
   Ldiff_UV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_0_out,
                 X => Ldiff_UV_del_1_0_IEEE);
Ldiff_UV_del_1_1_IEEE <= Ldiff_UV_del_1_1;
   Ldiff_UV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_1_out,
                 X => Ldiff_UV_del_1_1_IEEE);
Ldiff_UV_del_1_2_IEEE <= Ldiff_UV_del_1_2;
   Ldiff_UV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_2_out,
                 X => Ldiff_UV_del_1_2_IEEE);
Ldiff_UV_del_1_3_IEEE <= Ldiff_UV_del_1_3;
   Ldiff_UV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_3_out,
                 X => Ldiff_UV_del_1_3_IEEE);
Ldiff_UW_del_1_0_IEEE <= Ldiff_UW_del_1_0;
   Ldiff_UW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_0_out,
                 X => Ldiff_UW_del_1_0_IEEE);
Ldiff_UW_del_1_1_IEEE <= Ldiff_UW_del_1_1;
   Ldiff_UW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_1_out,
                 X => Ldiff_UW_del_1_1_IEEE);
Ldiff_UW_del_1_2_IEEE <= Ldiff_UW_del_1_2;
   Ldiff_UW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_2_out,
                 X => Ldiff_UW_del_1_2_IEEE);
Ldiff_UW_del_1_3_IEEE <= Ldiff_UW_del_1_3;
   Ldiff_UW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_3_out,
                 X => Ldiff_UW_del_1_3_IEEE);
Ldiff_VU_del_1_0_IEEE <= Ldiff_VU_del_1_0;
   Ldiff_VU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_0_out,
                 X => Ldiff_VU_del_1_0_IEEE);
Ldiff_VU_del_1_1_IEEE <= Ldiff_VU_del_1_1;
   Ldiff_VU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_1_out,
                 X => Ldiff_VU_del_1_1_IEEE);
Ldiff_VU_del_1_2_IEEE <= Ldiff_VU_del_1_2;
   Ldiff_VU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_2_out,
                 X => Ldiff_VU_del_1_2_IEEE);
Ldiff_VU_del_1_3_IEEE <= Ldiff_VU_del_1_3;
   Ldiff_VU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_3_out,
                 X => Ldiff_VU_del_1_3_IEEE);
Ldiff_VV_del_1_0_IEEE <= Ldiff_VV_del_1_0;
   Ldiff_VV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_0_out,
                 X => Ldiff_VV_del_1_0_IEEE);
Ldiff_VV_del_1_1_IEEE <= Ldiff_VV_del_1_1;
   Ldiff_VV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_1_out,
                 X => Ldiff_VV_del_1_1_IEEE);
Ldiff_VV_del_1_2_IEEE <= Ldiff_VV_del_1_2;
   Ldiff_VV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_2_out,
                 X => Ldiff_VV_del_1_2_IEEE);
Ldiff_VV_del_1_3_IEEE <= Ldiff_VV_del_1_3;
   Ldiff_VV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_3_out,
                 X => Ldiff_VV_del_1_3_IEEE);
Ldiff_VW_del_1_0_IEEE <= Ldiff_VW_del_1_0;
   Ldiff_VW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_0_out,
                 X => Ldiff_VW_del_1_0_IEEE);
Ldiff_VW_del_1_1_IEEE <= Ldiff_VW_del_1_1;
   Ldiff_VW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_1_out,
                 X => Ldiff_VW_del_1_1_IEEE);
Ldiff_VW_del_1_2_IEEE <= Ldiff_VW_del_1_2;
   Ldiff_VW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_2_out,
                 X => Ldiff_VW_del_1_2_IEEE);
Ldiff_VW_del_1_3_IEEE <= Ldiff_VW_del_1_3;
   Ldiff_VW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_3_out,
                 X => Ldiff_VW_del_1_3_IEEE);
Ldiff_WU_del_1_0_IEEE <= Ldiff_WU_del_1_0;
   Ldiff_WU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_0_out,
                 X => Ldiff_WU_del_1_0_IEEE);
Ldiff_WU_del_1_1_IEEE <= Ldiff_WU_del_1_1;
   Ldiff_WU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_1_out,
                 X => Ldiff_WU_del_1_1_IEEE);
Ldiff_WU_del_1_2_IEEE <= Ldiff_WU_del_1_2;
   Ldiff_WU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_2_out,
                 X => Ldiff_WU_del_1_2_IEEE);
Ldiff_WU_del_1_3_IEEE <= Ldiff_WU_del_1_3;
   Ldiff_WU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_3_out,
                 X => Ldiff_WU_del_1_3_IEEE);
Ldiff_WV_del_1_0_IEEE <= Ldiff_WV_del_1_0;
   Ldiff_WV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_0_out,
                 X => Ldiff_WV_del_1_0_IEEE);
Ldiff_WV_del_1_1_IEEE <= Ldiff_WV_del_1_1;
   Ldiff_WV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_1_out,
                 X => Ldiff_WV_del_1_1_IEEE);
Ldiff_WV_del_1_2_IEEE <= Ldiff_WV_del_1_2;
   Ldiff_WV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_2_out,
                 X => Ldiff_WV_del_1_2_IEEE);
Ldiff_WV_del_1_3_IEEE <= Ldiff_WV_del_1_3;
   Ldiff_WV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_3_out,
                 X => Ldiff_WV_del_1_3_IEEE);
Ldiff_WW_del_1_0_IEEE <= Ldiff_WW_del_1_0;
   Ldiff_WW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_0_out,
                 X => Ldiff_WW_del_1_0_IEEE);
Ldiff_WW_del_1_1_IEEE <= Ldiff_WW_del_1_1;
   Ldiff_WW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_1_out,
                 X => Ldiff_WW_del_1_1_IEEE);
Ldiff_WW_del_1_2_IEEE <= Ldiff_WW_del_1_2;
   Ldiff_WW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_2_out,
                 X => Ldiff_WW_del_1_2_IEEE);
Ldiff_WW_del_1_3_IEEE <= Ldiff_WW_del_1_3;
   Ldiff_WW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_3_out,
                 X => Ldiff_WW_del_1_3_IEEE);
R_U_0_IEEE <= R_U_0;
   R_U_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_0_out,
                 X => R_U_0_IEEE);
R_U_1_IEEE <= R_U_1;
   R_U_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_1_out,
                 X => R_U_1_IEEE);
R_U_2_IEEE <= R_U_2;
   R_U_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_2_out,
                 X => R_U_2_IEEE);
R_U_3_IEEE <= R_U_3;
   R_U_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_3_out,
                 X => R_U_3_IEEE);
R_V_0_IEEE <= R_V_0;
   R_V_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_0_out,
                 X => R_V_0_IEEE);
R_V_1_IEEE <= R_V_1;
   R_V_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_1_out,
                 X => R_V_1_IEEE);
R_V_2_IEEE <= R_V_2;
   R_V_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_2_out,
                 X => R_V_2_IEEE);
R_V_3_IEEE <= R_V_3;
   R_V_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_3_out,
                 X => R_V_3_IEEE);
R_W_0_IEEE <= R_W_0;
   R_W_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_0_out,
                 X => R_W_0_IEEE);
R_W_1_IEEE <= R_W_1;
   R_W_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_1_out,
                 X => R_W_1_IEEE);
R_W_2_IEEE <= R_W_2;
   R_W_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_2_out,
                 X => R_W_2_IEEE);
R_W_3_IEEE <= R_W_3;
   R_W_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_3_out,
                 X => R_W_3_IEEE);

Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_0_impl_out,
                 X => Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast);

Delay79No_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast <= Delay79No_out;
SharedReg943_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg235_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg235_out;
SharedReg44_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg933_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg933_out;
SharedReg927_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg227_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg227_out;
SharedReg335_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg937_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg298_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg298_out;
SharedReg299_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg299_out;
SharedReg222_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg222_out;
   MUX_Product108_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay79No_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg298_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg299_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg222_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg235_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg933_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg227_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg697_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg697_out;
SharedReg943_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg969_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg969_out;
SharedReg77_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg77_out;
SharedReg933_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg933_out;
SharedReg589_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg589_out;
SharedReg688_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg688_out;
SharedReg193_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg193_out;
SharedReg937_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg952_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg952_out;
SharedReg648_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg648_out;
SharedReg5_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg5_out;
   MUX_Product108_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg697_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg952_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg648_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg969_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg933_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg589_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg688_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg193_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product108_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_1_impl_out,
                 X => Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast);

SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg553_out;
SharedReg601_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg601_out;
SharedReg339_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg339_out;
SharedReg342_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg342_out;
SharedReg931_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg46_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg46_out;
SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg112_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg112_out;
SharedReg938_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg406_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg406_out;
SharedReg4_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg599_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg599_out;
   MUX_Product108_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg553_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg601_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg406_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg599_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg339_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg342_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg46_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg112_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg942_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg942_out;
SharedReg650_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg650_out;
SharedReg944_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg944_out;
SharedReg945_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg931_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg590_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg590_out;
SharedReg154_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg154_out;
SharedReg645_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg645_out;
SharedReg187_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg187_out;
SharedReg938_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg976_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg976_out;
SharedReg76_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg76_out;
SharedReg116_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg116_out;
   MUX_Product108_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg942_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg650_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg976_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg76_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg116_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg944_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg590_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg154_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg645_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg187_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product108_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_2_impl_out,
                 X => Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast);

SharedReg682_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg682_out;
SharedReg318_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg318_out;
SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg56_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg56_out;
SharedReg927_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg932_out;
SharedReg358_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg358_out;
SharedReg801_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg801_out;
SharedReg126_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg126_out;
SharedReg11_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg689_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg689_out;
SharedReg463_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg463_out;
SharedReg942_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg942_out;
   MUX_Product108_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg682_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg689_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg463_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg942_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg932_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg358_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg801_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg126_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg123_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg998_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg92_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg654_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg654_out;
SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg932_out;
SharedReg754_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg754_out;
SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg200_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg200_out;
SharedReg161_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg161_out;
SharedReg201_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg201_out;
SharedReg665_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg665_out;
SharedReg942_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg942_out;
   MUX_Product108_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg201_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg665_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg942_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg654_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg932_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg754_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg200_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg161_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product108_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_3_impl_out,
                 X => Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast);

SharedReg466_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg466_out;
SharedReg931_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg636_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg636_out;
SharedReg26_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg554_out;
SharedReg938_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg256_out;
SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg60_out;
SharedReg665_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg665_out;
SharedReg940_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product108_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg466_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg60_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg665_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg636_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg554_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_3_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_0_out,
                 Y => Delay1No6_out);

SharedReg675_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg675_out;
SharedReg931_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg758_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg758_out;
SharedReg172_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg172_out;
SharedReg708_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg708_out;
SharedReg935_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg666_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg666_out;
SharedReg947_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg947_out;
SharedReg938_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg138_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg138_out;
SharedReg664_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg664_out;
SharedReg749_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg749_out;
SharedReg940_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product108_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg675_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg664_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg749_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg758_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg708_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg666_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg947_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg138_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_3_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product110_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_0_impl_out,
                 X => Delay1No8_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast);

SharedReg225_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg943_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg338_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg226_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg226_out;
SharedReg372_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg372_out;
SharedReg927_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg301_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg301_out;
SharedReg936_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg234_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg234_out;
SharedReg264_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg264_out;
SharedReg940_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg941_out;
   MUX_Product110_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg264_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg338_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg226_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg372_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg301_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg936_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg234_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_0_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_0_out,
                 Y => Delay1No8_out);

SharedReg117_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg943_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
Delay90No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast <= Delay90No_out;
SharedReg958_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg958_out;
Delay94No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast <= Delay94No3_out;
SharedReg738_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg738_out;
SharedReg47_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg47_out;
SharedReg936_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg951_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg951_out;
SharedReg194_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg194_out;
SharedReg940_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg941_out;
   MUX_Product110_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg194_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay90No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg958_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay94No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg738_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg47_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg936_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg951_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_0_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product110_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_1_impl_out,
                 X => Delay1No10_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg600_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg600_out;
SharedReg330_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg330_out;
Delay1No217_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast <= Delay1No217_out;
SharedReg373_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg373_out;
SharedReg49_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg49_out;
SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg275_out;
SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg580_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg580_out;
SharedReg370_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg370_out;
SharedReg607_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg607_out;
SharedReg798_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg798_out;
SharedReg413_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg413_out;
   MUX_Product110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg600_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg330_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg607_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg798_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg413_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay1No217_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg373_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg49_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg580_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg370_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_1_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_0_out,
                 Y => Delay1No10_out);

SharedReg649_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg649_out;
SharedReg956_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg956_out;
SharedReg931_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg958_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg958_out;
SharedReg83_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg597_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg597_out;
SharedReg983_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg983_out;
SharedReg642_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg642_out;
SharedReg963_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg963_out;
SharedReg81_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg81_out;
SharedReg119_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg119_out;
SharedReg953_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg953_out;
SharedReg998_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg998_out;
   MUX_Product110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg649_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg956_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg119_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg953_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg998_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg958_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg597_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg983_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg642_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg963_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg81_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_1_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product110_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_2_impl_out,
                 X => Delay1No12_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg52_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
Delay94No6_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast <= Delay94No6_out;
SharedReg933_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg927_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg449_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg449_out;
Delay82No7_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast <= Delay82No7_out;
SharedReg90_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg90_out;
SharedReg851_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg851_out;
SharedReg694_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg694_out;
SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg561_out;
SharedReg846_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg846_out;
SharedReg248_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg248_out;
   MUX_Product110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg561_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg846_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg248_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay94No6_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg449_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay82No7_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg90_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg851_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg694_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_2_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_0_out,
                 Y => Delay1No12_out);

SharedReg700_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg954_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg954_out;
SharedReg637_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg637_out;
SharedReg933_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg705_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg705_out;
SharedReg54_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg99_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg99_out;
SharedReg658_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg658_out;
SharedReg983_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg983_out;
SharedReg709_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg709_out;
SharedReg1006_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1006_out;
SharedReg134_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg134_out;
Delay90No1_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast <= Delay90No1_out;
   MUX_Product110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg954_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1006_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg134_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay90No1_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg637_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg705_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg54_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg99_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg658_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg983_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg709_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_2_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product110_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_3_impl_out,
                 X => Delay1No14_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg545_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg545_out;
SharedReg465_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg465_out;
SharedReg550_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg550_out;
SharedReg626_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg626_out;
SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg937_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg208_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg208_out;
SharedReg941_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg796_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg796_out;
   MUX_Product110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg545_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg465_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg208_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg796_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg550_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg626_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg937_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_3_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_0_out,
                 Y => Delay1No14_out);

SharedReg979_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg979_out;
SharedReg211_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg1002_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1002_out;
SharedReg135_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg135_out;
SharedReg700_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg700_out;
SharedReg935_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg622_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg622_out;
SharedReg937_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg133_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg133_out;
SharedReg941_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg679_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg679_out;
   MUX_Product110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg979_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg133_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg679_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1002_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg135_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg700_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg622_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg937_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_3_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product109_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_0_impl_out,
                 X => Delay1No16_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg943_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg932_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg932_out;
SharedReg262_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg927_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg409_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg409_out;
Delay90No3_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast <= Delay90No3_out;
SharedReg296_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg296_out;
SharedReg938_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
Delay76No2_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast <= Delay76No2_out;
SharedReg490_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg490_out;
   MUX_Product109_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay76No2_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg490_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg932_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg409_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay90No3_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg296_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_0_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_0_out,
                 Y => Delay1No16_out);

SharedReg115_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg943_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg932_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg932_out;
SharedReg118_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg118_out;
SharedReg592_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg592_out;
SharedReg158_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg158_out;
SharedReg82_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg82_out;
SharedReg40_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg40_out;
SharedReg938_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg48_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg48_out;
Delay87No_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast <= Delay87No_out;
   MUX_Product109_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay87No_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg932_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg118_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg592_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg158_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg82_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg40_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_0_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product109_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_1_impl_out,
                 X => Delay1No18_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast);

SharedReg600_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg600_out;
SharedReg237_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg237_out;
Delay1No221_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast <= Delay1No221_out;
SharedReg519_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg519_out;
SharedReg931_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg231_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg486_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg486_out;
SharedReg74_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg74_out;
SharedReg272_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg272_out;
SharedReg411_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg411_out;
SharedReg524_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg524_out;
   MUX_Product109_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg600_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg272_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg411_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg524_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay1No221_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg519_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg486_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg74_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_1_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_0_out,
                 Y => Delay1No18_out);

SharedReg190_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg190_out;
SharedReg979_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg979_out;
SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg945_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg593_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg593_out;
SharedReg948_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg948_out;
SharedReg690_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg690_out;
SharedReg950_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg950_out;
SharedReg188_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg965_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg965_out;
SharedReg953_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg953_out;
SharedReg967_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg967_out;
   MUX_Product109_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg190_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg979_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg965_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg953_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg967_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg593_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg948_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg690_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg950_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_1_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product109_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_2_impl_out,
                 X => Delay1No20_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast);

SharedReg52_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg291_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg290_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg290_out;
SharedReg927_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg561_out;
SharedReg671_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg671_out;
SharedReg122_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg122_out;
SharedReg312_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg312_out;
SharedReg776_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
Delay97No1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast <= Delay97No1_out;
SharedReg941_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg941_out;
Delay68No4_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast <= Delay68No4_out;
   MUX_Product109_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay97No1_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay68No4_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg291_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg290_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg561_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg671_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg122_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg312_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_2_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_0_out,
                 Y => Delay1No20_out);

SharedReg700_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg988_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg988_out;
SharedReg681_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg681_out;
SharedReg98_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg617_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg617_out;
SharedReg661_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg174_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg174_out;
SharedReg160_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg160_out;
SharedReg948_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg948_out;
SharedReg962_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg962_out;
Delay100No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast <= Delay100No2_out;
SharedReg941_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg1009_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1009_out;
   MUX_Product109_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg988_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay100No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1009_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg681_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg617_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg661_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg174_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg160_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg948_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg962_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_2_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product109_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_3_impl_out,
                 X => Delay1No22_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast);

SharedReg475_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg475_out;
SharedReg25_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg625_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg625_out;
SharedReg175_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg175_out;
SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg782_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg782_out;
SharedReg938_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg427_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg427_out;
SharedReg420_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg420_out;
SharedReg462_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg462_out;
SharedReg526_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg526_out;
   MUX_Product109_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg475_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg420_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg462_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg526_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg625_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg175_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg782_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg427_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_3_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_0_out,
                 Y => Delay1No22_out);

SharedReg956_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg956_out;
SharedReg751_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg751_out;
SharedReg668_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg668_out;
SharedReg676_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg676_out;
SharedReg652_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg652_out;
SharedReg935_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg716_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg716_out;
SharedReg205_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg205_out;
SharedReg938_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
Delay100No4_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast <= Delay100No4_out;
SharedReg953_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg953_out;
SharedReg941_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg921_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg921_out;
   MUX_Product109_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg956_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg751_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg953_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg921_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg668_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg676_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg652_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg716_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg205_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay100No4_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_3_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_1_out,
                 Y => Delay1No23_out);

Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast <= Delay1No24_out;
Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast <= Delay1No25_out;
   Product111_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_0_impl_out,
                 X => Delay1No24_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No25_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast);

SharedReg79_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg943_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg363_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg363_out;
SharedReg932_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg932_out;
SharedReg8_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg927_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg935_out;
SharedReg232_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg232_out;
SharedReg408_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg408_out;
SharedReg296_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg296_out;
SharedReg939_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg442_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg442_out;
SharedReg941_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg941_out;
   MUX_Product111_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg442_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg363_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg932_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg935_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg232_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg408_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg296_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_0_impl_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_0_out,
                 Y => Delay1No24_out);

SharedReg692_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg692_out;
SharedReg943_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg641_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg641_out;
SharedReg932_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg932_out;
SharedReg153_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg153_out;
SharedReg737_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg737_out;
SharedReg935_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg935_out;
SharedReg962_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg962_out;
SharedReg80_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg80_out;
SharedReg113_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg113_out;
SharedReg939_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg691_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg691_out;
SharedReg941_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg941_out;
   MUX_Product111_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg692_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg691_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg641_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg932_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg153_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg737_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg935_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg962_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg80_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg113_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_0_impl_1_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_1_out,
                 Y => Delay1No25_out);

Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No26_out;
Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No27_out;
   Product111_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_1_impl_out,
                 X => Delay1No26_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No27_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg573_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg573_out;
Delay12No12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast <= Delay12No12_out;
SharedReg283_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg283_out;
SharedReg766_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg766_out;
SharedReg931_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg417_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg417_out;
SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg40_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg40_out;
SharedReg41_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg41_out;
SharedReg307_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg307_out;
SharedReg682_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg682_out;
SharedReg306_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg306_out;
   MUX_Product111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg573_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay12No12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg307_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg682_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg306_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg283_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg766_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg417_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg40_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg41_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_1_impl_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_0_out,
                 Y => Delay1No26_out);

SharedReg942_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg942_out;
SharedReg943_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg955_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg955_out;
Delay94No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast <= Delay94No1_out;
SharedReg931_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg732_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg732_out;
SharedReg698_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg698_out;
SharedReg605_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg605_out;
SharedReg150_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg150_out;
SharedReg188_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg976_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg976_out;
SharedReg638_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg638_out;
SharedReg967_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg967_out;
   MUX_Product111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg942_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg976_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg638_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg967_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg955_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay94No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg732_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg698_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg605_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg150_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_1_impl_1_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_1_out,
                 Y => Delay1No27_out);

Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No28_out;
Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No29_out;
   Product111_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_2_impl_out,
                 X => Delay1No28_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No29_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg163_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg163_out;
SharedReg387_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg387_out;
SharedReg932_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg933_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg927_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg848_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg848_out;
SharedReg754_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg754_out;
SharedReg246_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg246_out;
SharedReg759_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg759_out;
SharedReg538_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg538_out;
SharedReg771_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg771_out;
SharedReg324_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg324_out;
SharedReg942_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg942_out;
   MUX_Product111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg163_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg387_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg771_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg324_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg942_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg754_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg246_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg759_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg538_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_2_impl_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_0_out,
                 Y => Delay1No28_out);

SharedReg700_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg977_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg977_out;
SharedReg932_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg933_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg711_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg711_out;
SharedReg88_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg88_out;
SharedReg97_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg97_out;
SharedReg960_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg960_out;
SharedReg948_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg948_out;
SharedReg993_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg993_out;
SharedReg60_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg60_out;
SharedReg633_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg633_out;
SharedReg942_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg942_out;
   MUX_Product111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg977_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg60_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg633_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg942_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg711_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg88_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg97_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg960_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg948_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg993_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_2_impl_1_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_1_out,
                 Y => Delay1No29_out);

Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast <= Delay1No30_out;
Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast <= Delay1No31_out;
   Product111_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_3_impl_out,
                 X => Delay1No30_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No31_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast);

SharedReg504_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg249_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg515_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg515_out;
SharedReg56_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg56_out;
SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
Delay93No6_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast <= Delay93No6_out;
SharedReg938_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg838_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg838_out;
SharedReg505_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg505_out;
SharedReg810_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg810_out;
   MUX_Product111_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg838_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg505_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg810_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg515_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay93No6_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_3_impl_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_0_out,
                 Y => Delay1No30_out);

SharedReg943_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg943_out;
SharedReg944_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg944_out;
SharedReg990_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg990_out;
SharedReg92_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg745_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg745_out;
SharedReg935_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg749_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg749_out;
Delay93No3_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast <= Delay93No3_out;
SharedReg938_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg953_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg953_out;
SharedReg941_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg665_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg665_out;
   MUX_Product111_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg943_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg944_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg953_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg665_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg990_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg745_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg749_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay93No3_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_3_impl_1_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_1_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Product210_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_0_impl_out,
                 X => Delay1No32_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast);

SharedReg303_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg303_out;
SharedReg302_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg302_out;
SharedReg931_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg931_out;
Delay85No2_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast <= Delay85No2_out;
SharedReg45_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg927_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg402_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg402_out;
SharedReg457_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg457_out;
SharedReg937_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
Delay92No_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast <= Delay92No_out;
   MUX_Product210_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg302_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay92No_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay85No2_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg402_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg457_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg942_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg942_out;
SharedReg613_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg613_out;
SharedReg931_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg931_out;
Delay71No6_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast <= Delay71No6_out;
SharedReg643_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg643_out;
SharedReg740_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg740_out;
SharedReg948_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg948_out;
SharedReg993_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg993_out;
SharedReg937_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg9_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg9_out;
   MUX_Product210_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg942_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg613_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg9_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg931_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay71No6_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg643_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg740_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg948_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg993_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Product210_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_1_impl_out,
                 X => Delay1No34_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast);

Delay58No1_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast <= Delay58No1_out;
SharedReg239_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg239_out;
SharedReg500_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg500_out;
SharedReg10_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg931_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg271_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg271_out;
SharedReg574_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg574_out;
SharedReg927_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg439_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg439_out;
SharedReg781_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg781_out;
SharedReg403_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg403_out;
SharedReg522_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg522_out;
SharedReg497_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg497_out;
   MUX_Product210_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay58No1_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg239_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg403_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg522_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg497_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg500_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg271_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg574_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg439_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg781_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg987_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg987_out;
SharedReg663_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg663_out;
Delay81No8_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast <= Delay81No8_out;
SharedReg121_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg121_out;
SharedReg931_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg972_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg972_out;
SharedReg55_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg55_out;
SharedReg641_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg641_out;
SharedReg937_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg965_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg965_out;
SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg951_out;
SharedReg954_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg954_out;
   MUX_Product210_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg987_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg663_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg965_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg954_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay81No8_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg121_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg972_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg55_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg641_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Product210_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_2_impl_out,
                 X => Delay1No36_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast);

SharedReg503_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg503_out;
SharedReg579_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg579_out;
SharedReg352_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg352_out;
SharedReg933_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg927_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg50_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg50_out;
SharedReg514_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg514_out;
SharedReg385_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg385_out;
SharedReg800_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg800_out;
SharedReg783_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg783_out;
SharedReg399_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg399_out;
SharedReg941_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg469_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg469_out;
   MUX_Product210_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg503_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg579_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg399_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg469_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg352_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg50_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg514_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg385_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg800_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg783_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg953_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg953_out;
SharedReg954_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg954_out;
SharedReg209_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg209_out;
SharedReg933_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg933_out;
Delay84No1_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast <= Delay84No1_out;
SharedReg195_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg195_out;
SharedReg984_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg984_out;
SharedReg947_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg947_out;
SharedReg948_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg948_out;
SharedReg949_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg949_out;
SharedReg176_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg176_out;
SharedReg941_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg942_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg942_out;
   MUX_Product210_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg953_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg954_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg176_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg942_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg209_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay84No1_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg984_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg947_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg948_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg949_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Product210_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_3_impl_out,
                 X => Delay1No38_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast);

SharedReg72_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg569_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg323_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg323_out;
Delay83No4_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast <= Delay83No4_out;
SharedReg27_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg27_out;
Delay101No_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast <= Delay101No_out;
SharedReg927_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg383_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg383_out;
SharedReg938_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg288_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg288_out;
SharedReg748_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg748_out;
SharedReg254_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg254_out;
SharedReg940_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product210_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg748_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg254_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg323_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay83No4_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay101No_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg383_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg288_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg108_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg108_out;
SharedReg989_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg989_out;
SharedReg970_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg970_out;
Delay93No1_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast <= Delay93No1_out;
SharedReg136_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg136_out;
Delay97No2_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast <= Delay97No2_out;
SharedReg634_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg634_out;
SharedReg137_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg137_out;
SharedReg938_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg952_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg952_out;
SharedReg664_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg664_out;
SharedReg954_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg954_out;
SharedReg940_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product210_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg108_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg989_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg664_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg954_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg970_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay93No1_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg136_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay97No2_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg634_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg137_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg952_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product310_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_0_impl_out,
                 X => Delay1No40_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast);

SharedReg609_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg640_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg640_out;
SharedReg266_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg266_out;
Delay95No_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast <= Delay95No_out;
SharedReg604_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg604_out;
SharedReg927_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg446_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg446_out;
SharedReg334_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg334_out;
SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg329_out;
SharedReg938_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
Delay79No5_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast <= Delay79No5_out;
   MUX_Product310_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg640_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay79No5_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg266_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay95No_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg604_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg446_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg334_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg329_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_0_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_0_out,
                 Y => Delay1No40_out);

SharedReg695_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg695_out;
SharedReg152_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg614_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg614_out;
Delay97No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast <= Delay97No3_out;
SharedReg693_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg693_out;
SharedReg729_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg729_out;
SharedReg192_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg192_out;
SharedReg1013_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1013_out;
SharedReg155_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg155_out;
SharedReg938_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg651_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg651_out;
   MUX_Product310_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg695_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg651_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg614_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay97No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg729_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg192_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1013_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg155_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_0_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product310_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_1_impl_out,
                 X => Delay1No42_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast);

SharedReg243_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg781_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg781_out;
SharedReg942_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg306_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg306_out;
SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg481_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg481_out;
SharedReg281_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg281_out;
SharedReg927_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg453_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg453_out;
SharedReg3_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg412_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg412_out;
Delay64No4_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast <= Delay64No4_out;
   MUX_Product310_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg781_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg412_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay64No4_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg306_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg481_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg281_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg453_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_1_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_0_out,
                 Y => Delay1No42_out);

SharedReg700_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg53_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg942_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg124_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg129_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg129_out;
SharedReg947_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg947_out;
SharedReg971_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg971_out;
SharedReg654_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg654_out;
SharedReg935_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg951_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg951_out;
SharedReg114_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg114_out;
SharedReg202_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg202_out;
SharedReg998_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg998_out;
   MUX_Product310_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg114_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg998_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg129_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg947_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg971_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg654_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg951_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_1_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Product310_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_2_impl_out,
                 X => Delay1No44_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast);

SharedReg652_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg391_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg932_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg96_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg96_out;
SharedReg927_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg786_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg786_out;
SharedReg474_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg474_out;
SharedReg800_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg586_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg586_out;
SharedReg393_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg393_out;
SharedReg133_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg133_out;
SharedReg244_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg244_out;
SharedReg547_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg547_out;
   MUX_Product310_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg133_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg244_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg547_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg96_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg786_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg474_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg586_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg393_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_2_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_0_out,
                 Y => Delay1No44_out);

SharedReg700_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg998_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg932_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg752_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg752_out;
SharedReg615_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg615_out;
SharedReg1010_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1010_out;
SharedReg949_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg949_out;
SharedReg972_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg972_out;
SharedReg964_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg964_out;
SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg952_out;
SharedReg169_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg169_out;
SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg999_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg999_out;
   MUX_Product310_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg169_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg999_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg752_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg615_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1010_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg949_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg972_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg964_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_2_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product310_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_3_impl_out,
                 X => Delay1No46_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast);

SharedReg836_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg836_out;
SharedReg587_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg587_out;
SharedReg30_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg249_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg249_out;
SharedReg934_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg293_out;
SharedReg927_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg1006_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1006_out;
SharedReg427_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg427_out;
SharedReg563_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg23_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg24_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg24_out;
SharedReg527_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg527_out;
   MUX_Product310_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg836_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg587_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg527_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg30_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg249_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1006_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg427_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_3_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_0_out,
                 Y => Delay1No46_out);

SharedReg68_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg980_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg980_out;
SharedReg139_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg144_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg144_out;
SharedReg934_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg29_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg674_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg674_out;
SharedReg1006_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1006_out;
SharedReg28_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg28_out;
SharedReg939_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg748_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg748_out;
SharedReg170_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg170_out;
SharedReg997_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg997_out;
   MUX_Product310_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg980_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg748_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg170_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg997_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg139_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg144_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg674_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1006_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg28_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_3_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product410_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_0_impl_out,
                 X => Delay1No48_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast);

SharedReg768_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg768_out;
SharedReg610_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg610_out;
SharedReg487_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg487_out;
SharedReg233_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg233_out;
SharedReg39_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg927_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg363_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg363_out;
SharedReg375_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg375_out;
SharedReg937_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg330_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg330_out;
SharedReg940_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg231_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg231_out;
   MUX_Product410_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg768_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg610_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg330_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg231_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg487_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg233_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg363_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg375_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_0_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_0_out,
                 Y => Delay1No48_out);

Delay103No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast <= Delay103No_out;
SharedReg191_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg957_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg957_out;
SharedReg958_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg958_out;
SharedReg73_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg607_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg607_out;
SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg2_out;
SharedReg974_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg974_out;
SharedReg937_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg965_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg965_out;
SharedReg940_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg941_out;
   MUX_Product410_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay103No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg965_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg957_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg958_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg607_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg974_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_0_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product410_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_1_impl_out,
                 X => Delay1No50_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast);

SharedReg785_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg785_out;
SharedReg941_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg942_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg943_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
Delay98No_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast <= Delay98No_out;
Delay99No1_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast <= Delay99No1_out;
SharedReg927_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg364_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg364_out;
SharedReg378_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg378_out;
SharedReg938_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg938_out;
SharedReg5_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg5_out;
   MUX_Product410_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg785_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg378_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg938_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay98No_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay99No1_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg364_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_1_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_0_out,
                 Y => Delay1No50_out);

SharedReg203_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg941_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg942_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg943_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
Delay107No_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast <= Delay107No_out;
Delay98No2_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast <= Delay98No2_out;
SharedReg647_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg647_out;
SharedReg935_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg951_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg951_out;
SharedReg952_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg952_out;
SharedReg938_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg938_out;
SharedReg683_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg683_out;
   MUX_Product410_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg952_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg938_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg683_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay107No_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay98No2_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg647_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg951_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_1_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product410_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_2_impl_out,
                 X => Delay1No52_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast);

SharedReg564_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg564_out;
SharedReg931_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg932_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg130_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg130_out;
SharedReg927_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg50_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg50_out;
SharedReg843_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg843_out;
SharedReg540_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg540_out;
SharedReg320_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg320_out;
SharedReg241_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg241_out;
SharedReg251_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg251_out;
SharedReg941_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg476_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg476_out;
   MUX_Product410_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg564_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg251_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg476_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg130_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg50_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg843_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg540_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg320_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg241_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_2_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_0_out,
                 Y => Delay1No52_out);

SharedReg956_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg956_out;
SharedReg931_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg932_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg204_out;
SharedReg741_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg741_out;
SharedReg195_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg195_out;
SharedReg1005_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1005_out;
SharedReg1011_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1011_out;
SharedReg951_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg939_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg987_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg987_out;
SharedReg941_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg968_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg968_out;
   MUX_Product410_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg956_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg987_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg968_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg741_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1005_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1011_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_2_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product410_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_3_impl_out,
                 X => Delay1No54_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg624_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg624_out;
SharedReg817_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg817_out;
SharedReg825_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg825_out;
Delay87No7_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast <= Delay87No7_out;
SharedReg63_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg63_out;
SharedReg927_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg349_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg349_out;
SharedReg58_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg58_out;
SharedReg59_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg59_out;
SharedReg938_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg435_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg435_out;
SharedReg940_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product410_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg624_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg435_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg817_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg825_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay87No7_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg63_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg349_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg58_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg59_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_3_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_3_impl_0_out,
                 Y => Delay1No54_out);

SharedReg941_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg751_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg751_out;
SharedReg956_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg956_out;
SharedReg186_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg186_out;
Delay86No6_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast <= Delay86No6_out;
SharedReg173_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg173_out;
SharedReg633_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg633_out;
SharedReg168_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg168_out;
SharedReg206_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg206_out;
SharedReg207_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg207_out;
SharedReg938_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg954_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg954_out;
SharedReg940_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product410_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg751_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg954_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg956_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg186_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay86No6_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg173_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg633_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg168_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg206_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg207_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_3_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_3_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product510_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_0_impl_out,
                 X => Delay1No56_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast);

SharedReg43_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg43_out;
SharedReg7_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg308_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg308_out;
SharedReg341_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg341_out;
SharedReg_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg927_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg484_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg484_out;
SharedReg270_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg270_out;
SharedReg937_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg114_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg114_out;
SharedReg940_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg441_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg441_out;
   MUX_Product510_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg43_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg114_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg441_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg308_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg341_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg484_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg270_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_0_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_0_out,
                 Y => Delay1No56_out);

SharedReg639_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg639_out;
SharedReg685_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg685_out;
SharedReg969_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg969_out;
SharedReg945_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg73_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg595_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg688_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg688_out;
SharedReg962_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg962_out;
SharedReg937_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg938_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg151_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg940_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg940_out;
SharedReg977_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg977_out;
   MUX_Product510_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg639_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg685_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg977_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg969_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg688_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg962_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_0_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product510_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_1_impl_out,
                 X => Delay1No58_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast);

SharedReg940_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg942_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg523_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg523_out;
SharedReg931_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg263_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg263_out;
Delay82No6_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast <= Delay82No6_out;
SharedReg927_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg238_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg238_out;
SharedReg42_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg42_out;
SharedReg317_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg317_out;
SharedReg449_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg449_out;
   MUX_Product510_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg42_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg317_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg449_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg523_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg263_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay82No6_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg238_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_1_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_0_out,
                 Y => Delay1No58_out);

SharedReg940_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg941_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg942_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg942_out;
SharedReg166_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg166_out;
SharedReg931_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg157_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg157_out;
Delay93No4_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast <= Delay93No4_out;
SharedReg703_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg703_out;
SharedReg935_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg995_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg995_out;
SharedReg189_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg189_out;
SharedReg951_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg951_out;
SharedReg13_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg13_out;
   MUX_Product510_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg189_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg951_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg942_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg166_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg157_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay93No4_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg703_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg995_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_1_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product510_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_2_impl_out,
                 X => Delay1No60_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast);

SharedReg502_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg502_out;
SharedReg931_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg421_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg421_out;
SharedReg92_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg927_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg289_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg289_out;
SharedReg167_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg167_out;
SharedReg687_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg687_out;
SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg504_out;
SharedReg939_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg23_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg428_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg428_out;
SharedReg940_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product510_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg502_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg428_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg421_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg289_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg167_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg687_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_2_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_0_out,
                 Y => Delay1No60_out);

SharedReg171_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg931_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg945_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg945_out;
SharedReg204_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg204_out;
SharedReg713_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg713_out;
SharedReg753_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg753_out;
SharedReg132_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg132_out;
SharedReg704_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg704_out;
SharedReg21_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg939_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg94_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg94_out;
Delay80No9_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast <= Delay80No9_out;
SharedReg940_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product510_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg94_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay80No9_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg945_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg204_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg713_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg753_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg704_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_2_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product510_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_3_impl_out,
                 X => Delay1No62_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast);

SharedReg572_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg572_out;
SharedReg392_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg855_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg855_out;
SharedReg931_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg627_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg323_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg323_out;
SharedReg927_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg362_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg510_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg510_out;
SharedReg207_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg207_out;
SharedReg938_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg350_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg350_out;
SharedReg103_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg103_out;
   MUX_Product510_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg572_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg350_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg103_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg855_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg323_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg510_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg207_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_3_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_3_impl_0_out,
                 Y => Delay1No62_out);

SharedReg726_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg726_out;
SharedReg944_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg944_out;
SharedReg956_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg956_out;
SharedReg931_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg210_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg210_out;
SharedReg973_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg973_out;
SharedReg669_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg669_out;
Delay108No1_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast <= Delay108No1_out;
SharedReg951_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg93_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg93_out;
SharedReg938_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg954_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg954_out;
SharedReg917_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg917_out;
   MUX_Product510_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg726_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg944_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg954_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg917_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg956_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg210_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg973_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg669_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay108No1_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg93_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_3_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_3_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product610_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_1_impl_out,
                 X => Delay1No64_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast);

SharedReg498_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg498_out;
SharedReg941_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg556_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg556_out;
SharedReg539_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg539_out;
SharedReg686_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg686_out;
SharedReg333_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg333_out;
Delay96No6_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast <= Delay96No6_out;
SharedReg927_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg156_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg156_out;
SharedReg189_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg189_out;
SharedReg12_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
SharedReg797_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg797_out;
   MUX_Product610_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg498_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg189_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg797_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg556_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg539_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg686_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg333_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay96No6_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg156_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_1_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_0_out,
                 Y => Delay1No64_out);

SharedReg696_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg696_out;
SharedReg941_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg656_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg656_out;
Delay80No1_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast <= Delay80No1_out;
SharedReg125_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg125_out;
SharedReg605_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg605_out;
Delay108No_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast <= Delay108No_out;
SharedReg684_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg684_out;
SharedReg935_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg646_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg646_out;
SharedReg75_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg75_out;
SharedReg84_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg84_out;
SharedReg196_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg196_out;
   MUX_Product610_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg696_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg75_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg196_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg656_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay80No1_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg125_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg605_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay108No_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg684_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg646_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_1_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product610_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_3_impl_out,
                 X => Delay1No66_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg795_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg795_out;
SharedReg821_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg821_out;
SharedReg788_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg788_out;
SharedReg437_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg437_out;
SharedReg628_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg628_out;
SharedReg927_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg386_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg386_out;
SharedReg321_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg321_out;
SharedReg22_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg22_out;
SharedReg938_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg822_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg822_out;
SharedReg725_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg725_out;
   MUX_Product610_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg795_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg822_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg725_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg821_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg788_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg437_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg628_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg386_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg321_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg22_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_3_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_0_out,
                 Y => Delay1No66_out);

SharedReg941_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg1001_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg69_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg69_out;
SharedReg105_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
SharedReg972_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg972_out;
SharedReg670_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg670_out;
SharedReg664_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg664_out;
SharedReg630_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg630_out;
SharedReg951_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg93_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg93_out;
SharedReg938_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg954_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg954_out;
SharedReg185_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg185_out;
   MUX_Product610_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg954_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg185_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg69_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg972_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg670_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg664_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg630_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg93_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_3_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product710_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_1_impl_out,
                 X => Delay1No68_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast);

SharedReg940_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg454_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg454_out;
SharedReg86_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg943_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg784_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg784_out;
Delay85No3_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast <= Delay85No3_out;
SharedReg802_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg802_out;
SharedReg927_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg305_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg305_out;
SharedReg304_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg304_out;
SharedReg520_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg520_out;
SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg939_out;
   MUX_Product710_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg454_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg304_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg520_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg86_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg784_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay85No3_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg802_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg305_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_1_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_0_out,
                 Y => Delay1No68_out);

SharedReg940_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg128_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg128_out;
SharedReg198_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg943_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg969_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg969_out;
Delay93No2_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast <= Delay93No2_out;
SharedReg1003_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1003_out;
SharedReg736_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg736_out;
SharedReg935_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg975_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg975_out;
SharedReg952_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg952_out;
SharedReg951_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg951_out;
SharedReg939_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg939_out;
   MUX_Product710_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg952_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg951_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg939_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg198_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg969_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay93No2_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1003_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg736_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg975_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_1_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product710_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_3_impl_out,
                 X => Delay1No70_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
Delay1No216_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast <= Delay1No216_out;
SharedReg943_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg510_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg510_out;
SharedReg430_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg430_out;
SharedReg527_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg527_out;
SharedReg927_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg57_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg57_out;
SharedReg250_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg250_out;
SharedReg937_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg820_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg820_out;
SharedReg841_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg841_out;
SharedReg940_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product710_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No216_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg820_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg841_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg510_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg430_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg57_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg250_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_3_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_0_out,
                 Y => Delay1No70_out);

SharedReg941_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg931_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg943_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg944_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg944_out;
SharedReg947_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg947_out;
SharedReg961_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg961_out;
SharedReg677_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg677_out;
SharedReg168_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg168_out;
SharedReg951_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg937_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg722_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg722_out;
SharedReg976_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg976_out;
SharedReg940_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product710_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg722_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg976_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg944_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg947_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg961_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg677_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg168_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_3_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product810_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_1_impl_out,
                 X => Delay1No72_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast);

SharedReg535_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg941_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg684_out;
SharedReg943_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg349_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg349_out;
SharedReg934_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
SharedReg244_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg244_out;
SharedReg927_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
SharedReg935_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg188_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg347_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg347_out;
SharedReg51_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg51_out;
SharedReg777_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg777_out;
   MUX_Product810_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg347_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg51_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg777_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg349_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg244_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_1_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_0_out,
                 Y => Delay1No72_out);

SharedReg707_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg707_out;
SharedReg941_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg654_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg654_out;
SharedReg943_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg944_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg944_out;
SharedReg934_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg934_out;
SharedReg959_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg959_out;
SharedReg646_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg646_out;
SharedReg935_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg113_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg113_out;
SharedReg1007_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1007_out;
SharedReg162_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg162_out;
SharedReg976_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg976_out;
   MUX_Product810_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg707_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1007_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg162_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg976_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg654_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg944_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg959_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg646_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg113_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_1_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product810_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_3_impl_out,
                 X => Delay1No74_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast);

SharedReg544_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg544_out;
Delay1No219_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast <= Delay1No219_out;
SharedReg529_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg529_out;
Delay90No2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast <= Delay90No2_out;
SharedReg359_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg359_out;
SharedReg20_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg927_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg630_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg630_out;
SharedReg477_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg477_out;
SharedReg937_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg678_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg678_out;
SharedReg939_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg865_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg865_out;
   MUX_Product810_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg544_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No219_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg678_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg865_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg529_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay90No2_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg359_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg630_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg477_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_3_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_0_out,
                 Y => Delay1No74_out);

SharedReg219_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg219_out;
SharedReg931_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg145_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg145_out;
Delay96No7_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast <= Delay96No7_out;
SharedReg991_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg991_out;
SharedReg131_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg131_out;
Delay12No15_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast <= Delay12No15_out;
SharedReg137_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg137_out;
SharedReg964_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg964_out;
SharedReg937_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg922_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg922_out;
SharedReg939_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product810_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg219_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg922_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg145_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay96No7_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg991_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg131_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay12No15_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg137_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg964_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_3_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product910_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_1_impl_out,
                 X => Delay1No76_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast);

SharedReg700_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg941_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg311_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg311_out;
SharedReg764_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg764_out;
SharedReg49_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg49_out;
SharedReg644_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg644_out;
SharedReg759_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg759_out;
SharedReg927_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg927_out;
Delay79No4_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast <= Delay79No4_out;
SharedReg845_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg845_out;
SharedReg482_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg482_out;
SharedReg560_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg560_out;
SharedReg577_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg577_out;
   MUX_Product910_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg482_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg560_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg577_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg311_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg764_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg49_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg644_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg759_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg927_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay79No4_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg845_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_1_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_0_out,
                 Y => Delay1No76_out);

SharedReg163_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg163_out;
SharedReg941_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg968_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg968_out;
SharedReg956_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg956_out;
SharedReg83_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg687_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg687_out;
SharedReg933_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg933_out;
SharedReg603_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg603_out;
SharedReg91_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg91_out;
SharedReg938_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg938_out;
SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg985_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg985_out;
SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg939_out;
   MUX_Product910_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg163_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg985_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg939_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg968_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg956_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg933_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg603_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg91_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg938_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_1_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product910_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_3_impl_out,
                 X => Delay1No78_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast);

SharedReg831_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg831_out;
Delay1No223_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast <= Delay1No223_out;
SharedReg513_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg513_out;
SharedReg931_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg627_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg510_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg510_out;
SharedReg927_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
Delay18No2_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast <= Delay18No2_out;
SharedReg289_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
SharedReg508_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg508_out;
SharedReg33_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg33_out;
SharedReg939_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg839_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg839_out;
   MUX_Product910_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg831_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No223_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg33_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg839_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg513_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg510_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay18No2_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg508_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_3_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_0_out,
                 Y => Delay1No78_out);

SharedReg37_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg718_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg718_out;
SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg210_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg210_out;
SharedReg948_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg948_out;
SharedReg635_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg635_out;
SharedReg672_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg672_out;
SharedReg951_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg923_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg923_out;
SharedReg180_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg180_out;
SharedReg939_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
   MUX_Product910_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg180_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg718_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg210_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg948_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg635_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg672_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg923_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_3_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_1_out,
                 Y => Delay1No79_out);
   Inv_11_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_0_IEEE,
                 X => Delay1No80_out);
Inv_11_0 <= Inv_11_0_IEEE;

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => Delay1No80_out);
   Inv_11_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_1_IEEE,
                 X => Delay1No81_out);
Inv_11_1 <= Inv_11_1_IEEE;

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => Delay1No81_out);
   Inv_11_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_2_IEEE,
                 X => Delay1No82_out);
Inv_11_2 <= Inv_11_2_IEEE;

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => Delay1No82_out);
   Inv_11_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_3_IEEE,
                 X => Delay1No83_out);
Inv_11_3 <= Inv_11_3_IEEE;

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay1No83_out);
   Inv_12_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_0_IEEE,
                 X => Delay1No84_out);
Inv_12_0 <= Inv_12_0_IEEE;

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => Delay1No84_out);
   Inv_12_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_1_IEEE,
                 X => Delay1No85_out);
Inv_12_1 <= Inv_12_1_IEEE;

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => Delay1No85_out);
   Inv_12_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_2_IEEE,
                 X => Delay1No86_out);
Inv_12_2 <= Inv_12_2_IEEE;

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => Delay1No86_out);
   Inv_12_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_3_IEEE,
                 X => Delay1No87_out);
Inv_12_3 <= Inv_12_3_IEEE;

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => Delay1No87_out);
   Inv_13_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_0_IEEE,
                 X => Delay1No88_out);
Inv_13_0 <= Inv_13_0_IEEE;

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => Delay1No88_out);
   Inv_13_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_1_IEEE,
                 X => Delay1No89_out);
Inv_13_1 <= Inv_13_1_IEEE;

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => Delay1No89_out);
   Inv_13_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_2_IEEE,
                 X => Delay1No90_out);
Inv_13_2 <= Inv_13_2_IEEE;

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => Delay1No90_out);
   Inv_13_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_3_IEEE,
                 X => Delay1No91_out);
Inv_13_3 <= Inv_13_3_IEEE;

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => Delay1No91_out);
   Inv_21_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_0_IEEE,
                 X => Delay1No92_out);
Inv_21_0 <= Inv_21_0_IEEE;

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => Delay1No92_out);
   Inv_21_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_1_IEEE,
                 X => Delay1No93_out);
Inv_21_1 <= Inv_21_1_IEEE;

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => Delay1No93_out);
   Inv_21_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_2_IEEE,
                 X => Delay1No94_out);
Inv_21_2 <= Inv_21_2_IEEE;

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => Delay1No94_out);
   Inv_21_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_3_IEEE,
                 X => Delay1No95_out);
Inv_21_3 <= Inv_21_3_IEEE;

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => Delay1No95_out);
   Inv_22_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_0_IEEE,
                 X => Delay1No96_out);
Inv_22_0 <= Inv_22_0_IEEE;

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => Delay1No96_out);
   Inv_22_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_1_IEEE,
                 X => Delay1No97_out);
Inv_22_1 <= Inv_22_1_IEEE;

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => Delay1No97_out);
   Inv_22_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_2_IEEE,
                 X => Delay1No98_out);
Inv_22_2 <= Inv_22_2_IEEE;

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => Delay1No98_out);
   Inv_22_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_3_IEEE,
                 X => Delay1No99_out);
Inv_22_3 <= Inv_22_3_IEEE;

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => Delay1No99_out);
   Inv_23_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_0_IEEE,
                 X => Delay1No100_out);
Inv_23_0 <= Inv_23_0_IEEE;

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => Delay1No100_out);
   Inv_23_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_1_IEEE,
                 X => Delay1No101_out);
Inv_23_1 <= Inv_23_1_IEEE;

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => Delay1No101_out);
   Inv_23_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_2_IEEE,
                 X => Delay1No102_out);
Inv_23_2 <= Inv_23_2_IEEE;

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => Delay1No102_out);
   Inv_23_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_3_IEEE,
                 X => Delay1No103_out);
Inv_23_3 <= Inv_23_3_IEEE;

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => Delay1No103_out);
   Inv_31_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_0_IEEE,
                 X => Delay1No104_out);
Inv_31_0 <= Inv_31_0_IEEE;

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => Delay1No104_out);
   Inv_31_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_1_IEEE,
                 X => Delay1No105_out);
Inv_31_1 <= Inv_31_1_IEEE;

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => Delay1No105_out);
   Inv_31_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_2_IEEE,
                 X => Delay1No106_out);
Inv_31_2 <= Inv_31_2_IEEE;

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay1No106_out);
   Inv_31_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_3_IEEE,
                 X => Delay1No107_out);
Inv_31_3 <= Inv_31_3_IEEE;

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => Delay1No107_out);
   Inv_32_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_0_IEEE,
                 X => Delay1No108_out);
Inv_32_0 <= Inv_32_0_IEEE;

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => Delay1No108_out);
   Inv_32_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_1_IEEE,
                 X => Delay1No109_out);
Inv_32_1 <= Inv_32_1_IEEE;

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => Delay1No109_out);
   Inv_32_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_2_IEEE,
                 X => Delay1No110_out);
Inv_32_2 <= Inv_32_2_IEEE;

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => Delay1No110_out);
   Inv_32_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_3_IEEE,
                 X => Delay1No111_out);
Inv_32_3 <= Inv_32_3_IEEE;

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => Delay1No111_out);
   Inv_33_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_0_IEEE,
                 X => Delay1No112_out);
Inv_33_0 <= Inv_33_0_IEEE;

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => Delay1No112_out);
   Inv_33_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_1_IEEE,
                 X => Delay1No113_out);
Inv_33_1 <= Inv_33_1_IEEE;

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => Delay1No113_out);
   Inv_33_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_2_IEEE,
                 X => Delay1No114_out);
Inv_33_2 <= Inv_33_2_IEEE;

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => Delay1No114_out);
   Inv_33_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_3_IEEE,
                 X => Delay1No115_out);
Inv_33_3 <= Inv_33_3_IEEE;

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => Delay1No115_out);
   Inv_41_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_0_IEEE,
                 X => Delay1No116_out);
Inv_41_0 <= Inv_41_0_IEEE;

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => Delay1No116_out);
   Inv_41_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_1_IEEE,
                 X => Delay1No117_out);
Inv_41_1 <= Inv_41_1_IEEE;

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => Delay1No117_out);
   Inv_41_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_2_IEEE,
                 X => Delay1No118_out);
Inv_41_2 <= Inv_41_2_IEEE;

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => Delay1No118_out);
   Inv_41_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_3_IEEE,
                 X => Delay1No119_out);
Inv_41_3 <= Inv_41_3_IEEE;

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => Delay1No119_out);
   Inv_42_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_0_IEEE,
                 X => Delay1No120_out);
Inv_42_0 <= Inv_42_0_IEEE;

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => Delay1No120_out);
   Inv_42_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_1_IEEE,
                 X => Delay1No121_out);
Inv_42_1 <= Inv_42_1_IEEE;

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => Delay1No121_out);
   Inv_42_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_2_IEEE,
                 X => Delay1No122_out);
Inv_42_2 <= Inv_42_2_IEEE;

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => Delay1No122_out);
   Inv_42_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_3_IEEE,
                 X => Delay1No123_out);
Inv_42_3 <= Inv_42_3_IEEE;

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => Delay1No123_out);
   Inv_43_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_0_IEEE,
                 X => Delay1No124_out);
Inv_43_0 <= Inv_43_0_IEEE;

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => Delay1No124_out);
   Inv_43_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_1_IEEE,
                 X => Delay1No125_out);
Inv_43_1 <= Inv_43_1_IEEE;

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => Delay1No125_out);
   Inv_43_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_2_IEEE,
                 X => Delay1No126_out);
Inv_43_2 <= Inv_43_2_IEEE;

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => Delay1No126_out);
   Inv_43_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_3_IEEE,
                 X => Delay1No127_out);
Inv_43_3 <= Inv_43_3_IEEE;

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Add30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_0_impl_out,
                 X => Delay1No128_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg267_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg267_out;
SharedReg269_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg269_out;
SharedReg276_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg367_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg367_out;
SharedReg260_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg260_out;
SharedReg337_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg337_out;
SharedReg368_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg368_out;
SharedReg402_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg402_out;
SharedReg376_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg376_out;
SharedReg365_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg365_out;
SharedReg488_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg488_out;
Delay78No1_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast <= Delay78No1_out;
SharedReg405_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg405_out;
   MUX_Add30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg267_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg269_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg488_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay78No1_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg405_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg276_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg367_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg260_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg337_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg368_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg402_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg376_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg365_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_0_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_0_out,
                 Y => Delay1No128_out);

SharedReg892_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg892_out;
SharedReg223_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg223_out;
Delay56No3_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast <= Delay56No3_out;
SharedReg891_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg891_out;
SharedReg258_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg258_out;
SharedReg489_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg489_out;
SharedReg897_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg897_out;
SharedReg404_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg404_out;
SharedReg481_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg481_out;
SharedReg890_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg890_out;
SharedReg728_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg728_out;
SharedReg331_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg331_out;
SharedReg898_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg898_out;
   MUX_Add30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg892_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg223_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg728_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg331_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg898_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay56No3_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg891_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg258_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg489_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg897_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg404_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg481_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg890_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_0_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_1_impl_out,
                 X => Delay1No130_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg557_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg300_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg412_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg412_out;
SharedReg524_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg524_out;
SharedReg485_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg485_out;
SharedReg366_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg366_out;
Delay16No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast <= Delay16No_out;
SharedReg555_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg555_out;
SharedReg767_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg767_out;
SharedReg223_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg223_out;
SharedReg414_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg414_out;
SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg532_out;
SharedReg381_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg381_out;
   MUX_Add30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg414_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg381_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg412_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg524_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg485_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg366_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay16No_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg555_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg767_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg223_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_1_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_0_out,
                 Y => Delay1No130_out);

SharedReg521_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg521_out;
SharedReg901_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg901_out;
SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg734_out;
SharedReg314_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg314_out;
SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg734_out;
SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg734_out;
SharedReg340_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg340_out;
SharedReg598_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg598_out;
SharedReg602_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg602_out;
SharedReg731_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg731_out;
SharedReg652_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg652_out;
Delay13No41_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast <= Delay13No41_out;
SharedReg887_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg887_out;
   MUX_Add30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg521_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg901_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg652_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay13No41_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg887_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg314_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg340_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg598_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg602_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg731_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_1_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_2_impl_out,
                 X => Delay1No132_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast);

SharedReg315_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg774_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg774_out;
SharedReg874_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg874_out;
SharedReg859_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg859_out;
SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg316_out;
SharedReg433_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg433_out;
SharedReg322_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg322_out;
SharedReg253_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg253_out;
SharedReg310_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg310_out;
SharedReg847_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg847_out;
Delay90No4_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast <= Delay90No4_out;
SharedReg527_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg527_out;
SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg316_out;
   MUX_Add30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg774_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay90No4_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg527_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg874_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg859_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg316_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg433_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg322_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg253_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg310_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg847_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_2_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_0_out,
                 Y => Delay1No132_out);

SharedReg914_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg914_out;
SharedReg325_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg325_out;
SharedReg911_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg911_out;
SharedReg527_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg527_out;
SharedReg503_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg503_out;
SharedReg479_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg479_out;
SharedReg741_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg741_out;
SharedReg509_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg509_out;
Delay68No3_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast <= Delay68No3_out;
SharedReg652_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg652_out;
SharedReg631_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg631_out;
SharedReg615_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg615_out;
SharedReg901_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg901_out;
   MUX_Add30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg914_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg325_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg631_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg615_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg901_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg911_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg527_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg503_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg479_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg741_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg509_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay68No3_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg652_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_2_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Add30_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_3_impl_out,
                 X => Delay1No134_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast);

SharedReg436_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg436_out;
SharedReg527_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg527_out;
SharedReg397_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg397_out;
Delay89No1_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast <= Delay89No1_out;
SharedReg568_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg287_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg287_out;
SharedReg787_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg787_out;
SharedReg582_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg582_out;
Delay7No_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast <= Delay7No_out;
SharedReg530_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg530_out;
SharedReg803_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg803_out;
SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg396_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg396_out;
   MUX_Add30_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg436_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg527_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg803_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg396_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg397_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay89No1_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg568_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg287_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg787_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg582_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay7No_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg530_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_3_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_0_out,
                 Y => Delay1No134_out);

SharedReg915_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg915_out;
SharedReg748_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg748_out;
SharedReg904_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg904_out;
SharedReg902_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg623_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg623_out;
SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg741_out;
SharedReg917_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg917_out;
SharedReg819_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg819_out;
SharedReg543_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg543_out;
SharedReg907_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg907_out;
SharedReg895_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg895_out;
SharedReg629_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg629_out;
SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg741_out;
   MUX_Add30_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg915_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg748_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg895_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg629_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg904_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg623_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg741_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg917_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg819_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg543_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg907_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_3_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Add110_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_1_impl_out,
                 X => Delay1No136_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg853_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg853_out;
SharedReg440_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg440_out;
SharedReg846_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg846_out;
SharedReg799_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg799_out;
Delay85No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast <= Delay85No4_out;
SharedReg345_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg345_out;
Delay3No2_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast <= Delay3No2_out;
SharedReg268_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg268_out;
SharedReg351_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg351_out;
SharedReg265_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg265_out;
SharedReg518_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg518_out;
Delay94No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast <= Delay94No4_out;
SharedReg349_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg349_out;
   MUX_Add110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg853_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg440_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg518_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay94No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg349_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg846_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay85No4_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg345_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay3No2_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg268_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg351_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg265_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_1_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_0_out,
                 Y => Delay1No136_out);

Delay89No2_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast <= Delay89No2_out;
SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg682_out;
SharedReg700_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg700_out;
SharedReg897_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg897_out;
Delay79No8_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast <= Delay79No8_out;
SharedReg899_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg899_out;
SharedReg268_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg268_out;
SharedReg734_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg734_out;
SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg682_out;
SharedReg886_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg886_out;
SharedReg896_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg896_out;
SharedReg889_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg889_out;
SharedReg761_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg761_out;
   MUX_Add110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay89No2_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg896_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg889_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg761_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg700_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg897_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay79No8_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg268_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg734_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg682_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg886_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_1_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Add110_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_2_impl_out,
                 X => Delay1No138_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg783_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg461_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg461_out;
SharedReg383_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg383_out;
SharedReg350_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg350_out;
SharedReg782_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg782_out;
Delay85No5_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast <= Delay85No5_out;
SharedReg395_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg395_out;
SharedReg241_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg241_out;
Delay6No9_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast <= Delay6No9_out;
SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg419_out;
SharedReg781_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg781_out;
SharedReg468_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg468_out;
SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg511_out;
   MUX_Add110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg461_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg781_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg468_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg511_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg383_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg350_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg782_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay85No5_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg395_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg241_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No9_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg419_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_2_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_0_out,
                 Y => Delay1No138_out);

SharedReg908_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg711_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg711_out;
SharedReg902_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg245_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg245_out;
SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg638_out;
SharedReg910_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg910_out;
SharedReg507_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg507_out;
SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg638_out;
SharedReg769_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg769_out;
SharedReg415_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg415_out;
SharedReg906_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg906_out;
SharedReg746_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg746_out;
SharedReg905_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg905_out;
   MUX_Add110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg711_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg906_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg746_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg905_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg902_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg245_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg910_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg507_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg638_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg769_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg415_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_2_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Add110_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_3_impl_out,
                 X => Delay1No140_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg516_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg516_out;
SharedReg567_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg567_out;
SharedReg806_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg806_out;
SharedReg882_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg882_out;
SharedReg878_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg878_out;
Delay4No7_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast <= Delay4No7_out;
Delay19No_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast <= Delay19No_out;
SharedReg837_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg837_out;
SharedReg361_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg361_out;
SharedReg581_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg581_out;
SharedReg814_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg814_out;
SharedReg826_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg826_out;
SharedReg789_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg789_out;
   MUX_Add110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg516_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg567_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg814_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg826_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg789_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg806_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg882_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg878_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No7_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay19No_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg837_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg361_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg581_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_3_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_0_out,
                 Y => Delay1No140_out);

SharedReg748_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg748_out;
SharedReg912_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg912_out;
SharedReg909_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg716_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg716_out;
SharedReg911_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg911_out;
SharedReg563_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg563_out;
SharedReg880_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg880_out;
SharedReg916_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg916_out;
Delay73No2_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast <= Delay73No2_out;
SharedReg817_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg817_out;
SharedReg548_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg548_out;
SharedReg913_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg913_out;
Delay87No8_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast <= Delay87No8_out;
   MUX_Add110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg748_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg912_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg548_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg913_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay87No8_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg909_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg716_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg911_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg563_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg880_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg916_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay73No2_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg817_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_3_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Add101_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_1_impl_out,
                 X => Delay1No142_out_to_Add101_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Add101_1_impl_parent_implementedSystem_port_1_cast);

SharedReg452_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg452_out;
SharedReg380_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg380_out;
SharedReg350_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg350_out;
SharedReg760_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg423_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg781_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg781_out;
Delay3No10_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast <= Delay3No10_out;
SharedReg573_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg573_out;
Delay6No_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast <= Delay6No_out;
SharedReg483_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg483_out;
SharedReg501_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg501_out;
SharedReg420_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg420_out;
SharedReg353_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg353_out;
   MUX_Add101_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg452_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg380_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg501_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg420_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg353_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg350_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg781_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay3No10_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg573_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg483_out_to_MUX_Add101_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_1_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_1_impl_0_out,
                 Y => Delay1No142_out);

SharedReg905_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg905_out;
SharedReg575_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg575_out;
SharedReg420_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg420_out;
SharedReg682_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg682_out;
SharedReg608_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg608_out;
SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg797_out;
SharedReg303_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg303_out;
SharedReg494_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg494_out;
SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg797_out;
SharedReg598_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg598_out;
SharedReg418_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg418_out;
SharedReg700_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg700_out;
SharedReg652_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg652_out;
   MUX_Add101_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg905_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg575_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg418_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg700_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg652_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg420_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg682_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg608_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg303_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg494_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg797_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg598_out_to_MUX_Add101_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_1_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_1_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add111_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_1_impl_out,
                 X => Delay1No144_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg763_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg763_out;
SharedReg536_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg536_out;
SharedReg504_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg504_out;
SharedReg434_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg434_out;
SharedReg765_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg765_out;
SharedReg778_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg778_out;
SharedReg573_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg573_out;
SharedReg780_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg780_out;
Delay6No4_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast <= Delay6No4_out;
SharedReg346_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg346_out;
SharedReg313_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg313_out;
SharedReg472_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg472_out;
SharedReg394_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg394_out;
   MUX_Add111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg763_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg536_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg313_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg472_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg394_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg504_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg434_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg765_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg778_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg573_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg780_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No4_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg346_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_1_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_0_out,
                 Y => Delay1No144_out);

SharedReg701_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg701_out;
SharedReg496_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg496_out;
SharedReg277_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg277_out;
SharedReg899_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg373_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg373_out;
SharedReg693_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg693_out;
SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg711_out;
SharedReg388_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg388_out;
SharedReg845_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg845_out;
SharedReg900_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg900_out;
SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg711_out;
SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg911_out;
SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg911_out;
   MUX_Add111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg701_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg496_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg911_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg277_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg373_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg693_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg711_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg388_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg845_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg900_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_1_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Add111_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_2_impl_out,
                 X => Delay1No146_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg360_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg360_out;
SharedReg384_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg384_out;
Delay77No2_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast <= Delay77No2_out;
SharedReg459_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg459_out;
SharedReg425_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg576_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg576_out;
SharedReg464_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg773_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg773_out;
SharedReg278_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg278_out;
SharedReg281_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg281_out;
SharedReg528_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg528_out;
SharedReg836_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg836_out;
Delay87No5_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_13_cast <= Delay87No5_out;
   MUX_Add111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg360_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg384_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg528_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg836_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay87No5_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay77No2_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg459_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg576_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg773_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg278_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg281_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_2_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_2_impl_0_out,
                 Y => Delay1No146_out);

SharedReg660_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg660_out;
SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg615_out;
SharedReg844_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg844_out;
SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg615_out;
SharedReg682_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg682_out;
SharedReg894_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg894_out;
SharedReg623_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg623_out;
SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg903_out;
SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg903_out;
SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg711_out;
SharedReg252_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg252_out;
SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg711_out;
SharedReg632_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg632_out;
   MUX_Add111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg660_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg252_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg632_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg844_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg615_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg682_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg894_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg623_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg903_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg711_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_2_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_2_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Add121_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_3_impl_out,
                 X => Delay1No148_out_to_Add121_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Add121_3_impl_parent_implementedSystem_port_1_cast);

Delay7No7_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast <= Delay7No7_out;
SharedReg289_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg289_out;
SharedReg792_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg792_out;
SharedReg582_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg582_out;
SharedReg825_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg825_out;
SharedReg791_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg791_out;
SharedReg883_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg883_out;
SharedReg928_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg928_out;
   MUX_Add121_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No7_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg289_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg792_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg582_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg825_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg791_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg883_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg928_out_to_MUX_Add121_3_impl_0_parent_implementedSystem_port_8_cast,
                 iSel => MUX_Add121_3_impl_0_LUT_out,
                 oMux => MUX_Add121_3_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_0_out,
                 Y => Delay1No148_out);

SharedReg673_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg326_out;
SharedReg808_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg808_out;
SharedReg830_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg830_out;
SharedReg748_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg748_out;
SharedReg716_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg716_out;
SharedReg866_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg866_out;
SharedReg880_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg880_out;
   MUX_Add121_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg808_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg830_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg748_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg716_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg866_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg880_out_to_MUX_Add121_3_impl_1_parent_implementedSystem_port_8_cast,
                 iSel => MUX_Add121_3_impl_1_LUT_out,
                 oMux => MUX_Add121_3_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_3_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Add141_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_0_impl_out,
                 X => Delay1No150_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast);

SharedReg297_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg443_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg443_out;
SharedReg444_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg444_out;
SharedReg537_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg537_out;
SharedReg447_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg447_out;
SharedReg229_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg229_out;
SharedReg236_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg236_out;
SharedReg224_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg224_out;
SharedReg274_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg274_out;
SharedReg369_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg369_out;
SharedReg303_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg303_out;
SharedReg451_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg451_out;
SharedReg402_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg402_out;
   MUX_Add141_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg443_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg303_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg451_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg402_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg444_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg537_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg447_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg229_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg236_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg224_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg274_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg369_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_0_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_0_out,
                 Y => Delay1No150_out);

SharedReg493_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg493_out;
SharedReg403_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg735_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg735_out;
SharedReg886_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg886_out;
SharedReg889_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg889_out;
SharedReg336_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg336_out;
Delay59No_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast <= Delay59No_out;
SharedReg257_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg257_out;
SharedReg727_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg727_out;
SharedReg591_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg591_out;
SharedReg344_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg344_out;
SharedReg893_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg893_out;
SharedReg598_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg598_out;
   MUX_Add141_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg493_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg344_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg893_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg598_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg735_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg886_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg889_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg336_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay59No_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg257_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg727_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg591_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_0_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Add141_1_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Add141_1_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Add141_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_1_impl_out,
                 X => Delay1No152_out_to_Add141_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Add141_1_impl_parent_implementedSystem_port_1_cast);

SharedReg491_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg491_out;
SharedReg261_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg261_out;
SharedReg532_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg532_out;
SharedReg779_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg779_out;
SharedReg439_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg439_out;
SharedReg522_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg522_out;
SharedReg343_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg343_out;
SharedReg379_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg379_out;
SharedReg762_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg762_out;
SharedReg371_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg371_out;
SharedReg273_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg273_out;
SharedReg775_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg775_out;
SharedReg455_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg455_out;
   MUX_Add141_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg491_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg261_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg273_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg775_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg455_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg532_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg779_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg439_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg522_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg343_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg379_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg762_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg371_out_to_MUX_Add141_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_1_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_1_impl_0_out,
                 Y => Delay1No152_out);

SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg727_out;
SharedReg892_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg892_out;
SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg727_out;
SharedReg704_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg704_out;
SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg888_out;
SharedReg332_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg332_out;
SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg638_out;
SharedReg643_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg643_out;
SharedReg852_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg852_out;
SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg888_out;
SharedReg598_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg598_out;
SharedReg899_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg899_out;
SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg638_out;
   MUX_Add141_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg892_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg598_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg899_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg727_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg704_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg332_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg638_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg643_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg852_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg888_out_to_MUX_Add141_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_1_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_1_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Add17_3_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Add17_3_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Add17_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add17_3_impl_out,
                 X => Delay1No154_out_to_Add17_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Add17_3_impl_parent_implementedSystem_port_1_cast);

SharedReg396_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg396_out;
SharedReg355_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg355_out;
SharedReg823_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg823_out;
SharedReg866_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg866_out;
SharedReg461_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg461_out;
SharedReg322_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg322_out;
SharedReg822_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg822_out;
SharedReg356_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg356_out;
SharedReg525_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg525_out;
SharedReg546_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg546_out;
SharedReg424_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg424_out;
SharedReg827_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg827_out;
Delay98No1_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_13_cast <= Delay98No1_out;
   MUX_Add17_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg396_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg355_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg424_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg827_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay98No1_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg823_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg866_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg461_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg322_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg822_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg356_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg525_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg546_out_to_MUX_Add17_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add17_3_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add17_3_impl_0_out,
                 Y => Delay1No154_out);

SharedReg741_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg741_out;
SharedReg664_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg664_out;
SharedReg816_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg816_out;
SharedReg911_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg911_out;
SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg744_out;
SharedReg615_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg615_out;
SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg744_out;
SharedReg652_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg652_out;
SharedReg711_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg711_out;
SharedReg390_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg390_out;
SharedReg467_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg467_out;
Delay48No_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_12_cast <= Delay48No_out;
SharedReg914_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg914_out;
   MUX_Add17_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg741_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg664_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg467_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay48No_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg914_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg816_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg911_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg615_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg744_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg652_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg711_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg390_out_to_MUX_Add17_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add17_3_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add17_3_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Add22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Add22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Add22_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add22_3_impl_out,
                 X => Delay1No156_out_to_Add22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Add22_3_impl_parent_implementedSystem_port_1_cast);

Delay4No9_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_1_cast <= Delay4No9_out;
SharedReg549_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg549_out;
SharedReg807_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg807_out;
SharedReg824_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg438_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg438_out;
SharedReg877_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg877_out;
SharedReg858_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg856_out;
SharedReg422_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg422_out;
SharedReg929_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg929_out;
SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg856_out;
   MUX_Add22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No9_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg549_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg807_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg438_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg877_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg856_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg422_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg929_out_to_MUX_Add22_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add22_3_impl_0_LUT_out,
                 oMux => MUX_Add22_3_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_3_impl_0_out,
                 Y => Delay1No156_out);

SharedReg757_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg757_out;
SharedReg755_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg755_out;
SharedReg826_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg826_out;
SharedReg818_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg818_out;
SharedReg879_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg879_out;
SharedReg912_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
SharedReg623_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg623_out;
SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg917_out;
SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg917_out;
SharedReg748_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg748_out;
SharedReg581_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg581_out;
   MUX_Add22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg757_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg755_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg581_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg826_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg818_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg879_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg623_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg917_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg748_out_to_MUX_Add22_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add22_3_impl_1_LUT_out,
                 oMux => MUX_Add22_3_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_3_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product112_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_1_impl_out,
                 X => Delay1No158_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast);

SharedReg700_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg499_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg499_out;
SharedReg159_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg159_out;
SharedReg850_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg850_out;
SharedReg420_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg420_out;
SharedReg934_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
SharedReg578_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg578_out;
SharedReg242_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg242_out;
SharedReg935_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg374_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg255_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg255_out;
SharedReg196_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg196_out;
   MUX_Product112_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg499_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg255_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg196_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg159_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg850_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg420_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg578_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg242_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product112_1_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_0_out,
                 Y => Delay1No158_out);

SharedReg652_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg19_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg120_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg979_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg979_out;
SharedReg944_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg944_out;
SharedReg934_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg934_out;
SharedReg946_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg946_out;
SharedReg947_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg947_out;
SharedReg935_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg975_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg975_out;
SharedReg85_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg85_out;
   MUX_Product112_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg975_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg85_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg979_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg944_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg946_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg947_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product112_1_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product112_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_2_impl_out,
                 X => Delay1No160_out_to_Product112_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product112_2_impl_parent_implementedSystem_port_1_cast);

SharedReg240_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg240_out;
SharedReg15_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg932_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg759_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg759_out;
Delay1No222_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast <= Delay1No222_out;
SharedReg279_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg279_out;
SharedReg284_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg284_out;
SharedReg934_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg934_out;
SharedReg458_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg458_out;
SharedReg533_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg533_out;
SharedReg799_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg799_out;
SharedReg941_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg431_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg431_out;
   MUX_Product112_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg240_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg799_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg431_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg759_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay1No222_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg279_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg284_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg934_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg458_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg533_out_to_MUX_Product112_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product112_2_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_0_out,
                 Y => Delay1No160_out);

SharedReg940_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg164_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg164_out;
SharedReg932_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg943_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg970_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg970_out;
SharedReg64_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg64_out;
SharedReg934_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg934_out;
SharedReg699_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg699_out;
SharedReg949_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg949_out;
SharedReg950_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg950_out;
SharedReg941_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg941_out;
SharedReg61_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg61_out;
   MUX_Product112_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg164_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg950_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg941_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg61_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg970_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg64_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg934_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg699_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg949_out_to_MUX_Product112_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product112_2_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_2_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product113_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_2_impl_out,
                 X => Delay1No162_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast);

SharedReg682_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg682_out;
SharedReg770_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg770_out;
SharedReg932_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg655_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg655_out;
SharedReg18_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
Delay96No3_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_7_cast <= Delay96No3_out;
Delay94No5_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_8_cast <= Delay94No5_out;
SharedReg577_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg577_out;
SharedReg936_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg17_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg17_out;
SharedReg772_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg772_out;
   MUX_Product113_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg682_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg770_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg17_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg772_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg655_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay96No3_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay94No5_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg577_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product113_2_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_2_impl_0_out,
                 Y => Delay1No162_out);

SharedReg197_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg197_out;
SharedReg683_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg683_out;
SharedReg932_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg87_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg87_out;
SharedReg657_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg657_out;
SharedReg149_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg149_out;
Delay108No2_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_7_cast <= Delay108No2_out;
Delay111No_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_8_cast <= Delay111No_out;
SharedReg948_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg948_out;
SharedReg936_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg127_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg127_out;
SharedReg952_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg952_out;
   MUX_Product113_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg197_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg683_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg127_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg952_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg87_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg657_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg149_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay108No2_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay111No_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg948_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product113_2_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_2_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product113_3_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product113_3_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product113_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_3_impl_out,
                 X => Delay1No164_out_to_Product113_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product113_3_impl_parent_implementedSystem_port_1_cast);

SharedReg107_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg942_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg942_out;
SharedReg812_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg812_out;
SharedReg31_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg31_out;
Delay96No4_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_5_cast <= Delay96No4_out;
SharedReg933_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg400_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg400_out;
SharedReg517_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg517_out;
SharedReg526_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg526_out;
SharedReg937_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg71_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg71_out;
SharedReg939_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
Delay54No_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_13_cast <= Delay54No_out;
   MUX_Product113_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg71_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay54No_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg812_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay96No4_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg517_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg526_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product113_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product113_3_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_3_impl_0_out,
                 Y => Delay1No164_out);

SharedReg221_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg942_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg942_out;
SharedReg1000_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1000_out;
SharedReg178_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg178_out;
Delay107No1_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_5_cast <= Delay107No1_out;
SharedReg933_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg933_out;
Delay97No_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_7_cast <= Delay97No_out;
SharedReg109_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg109_out;
SharedReg951_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg937_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg722_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg722_out;
SharedReg939_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg1008_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1008_out;
   MUX_Product113_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg722_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1008_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1000_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay107No1_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay97No_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg109_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product113_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product113_3_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_3_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product103_2_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product103_2_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product103_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product103_2_impl_out,
                 X => Delay1No166_out_to_Product103_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product103_2_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg495_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg495_out;
SharedReg932_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg199_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg199_out;
Delay1No215_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_5_cast <= Delay1No215_out;
SharedReg687_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg687_out;
SharedReg506_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg506_out;
SharedReg533_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg533_out;
SharedReg935_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg935_out;
Delay93No5_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_10_cast <= Delay93No5_out;
SharedReg937_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg784_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg784_out;
SharedReg13_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg13_out;
   MUX_Product103_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg495_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg784_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg199_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay1No215_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg506_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg533_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay93No5_out_to_MUX_Product103_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product103_2_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product103_2_impl_0_out,
                 Y => Delay1No166_out);

SharedReg652_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg701_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg701_out;
SharedReg932_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg124_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg124_out;
SharedReg931_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg78_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg78_out;
SharedReg949_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg949_out;
SharedReg165_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg935_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg935_out;
Delay100No1_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_10_cast <= Delay100No1_out;
SharedReg937_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg964_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg964_out;
SharedReg85_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg85_out;
   MUX_Product103_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg701_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg964_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg85_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg78_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg949_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg935_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay100No1_out_to_MUX_Product103_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product103_2_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product103_2_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product103_3_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product103_3_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product103_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product103_3_impl_out,
                 X => Delay1No168_out_to_Product103_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product103_3_impl_parent_implementedSystem_port_1_cast);

SharedReg717_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg717_out;
SharedReg815_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg815_out;
SharedReg65_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg668_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg668_out;
Delay79No7_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_5_cast <= Delay79No7_out;
SharedReg933_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg842_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg842_out;
Delay84No4_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_8_cast <= Delay84No4_out;
SharedReg936_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg936_out;
Delay87No6_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_10_cast <= Delay87No6_out;
SharedReg790_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg790_out;
SharedReg939_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg861_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg861_out;
   MUX_Product103_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg717_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg815_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg790_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg861_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg668_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay79No7_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg842_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay84No4_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg936_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay87No6_out_to_MUX_Product103_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product103_3_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product103_3_impl_0_out,
                 Y => Delay1No168_out);

SharedReg918_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
Delay87No3_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_2_cast <= Delay87No3_out;
SharedReg177_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg177_out;
SharedReg146_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg146_out;
SharedReg1010_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1010_out;
SharedReg933_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg670_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg670_out;
SharedReg110_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg110_out;
SharedReg936_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg936_out;
Delay96No2_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_10_cast <= Delay96No2_out;
SharedReg964_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg964_out;
SharedReg939_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg953_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg953_out;
   MUX_Product103_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay87No3_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg964_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg953_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg177_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg146_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1010_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg670_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg110_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg936_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay96No2_out_to_MUX_Product103_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product103_3_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product103_3_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product106_3_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product106_3_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product106_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product106_3_impl_out,
                 X => Delay1No170_out_to_Product106_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product106_3_impl_parent_implementedSystem_port_1_cast);

SharedReg584_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg584_out;
SharedReg942_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg942_out;
SharedReg943_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg793_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg793_out;
SharedReg355_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg355_out;
SharedReg933_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg794_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg429_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg429_out;
SharedReg356_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg356_out;
SharedReg585_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg585_out;
SharedReg71_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg71_out;
Delay75No1_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_12_cast <= Delay75No1_out;
SharedReg840_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg840_out;
   MUX_Product106_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg584_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg71_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay75No1_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg840_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg793_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg355_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg429_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg356_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg585_out_to_MUX_Product106_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product106_3_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product106_3_impl_0_out,
                 Y => Delay1No170_out);

SharedReg918_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg942_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg942_out;
SharedReg943_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg980_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg980_out;
SharedReg947_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg947_out;
SharedReg933_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg184_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg184_out;
SharedReg935_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg935_out;
SharedReg938_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg36_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg36_out;
SharedReg722_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg722_out;
SharedReg148_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg148_out;
SharedReg966_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg966_out;
   MUX_Product106_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg722_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg148_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg966_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg980_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg947_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg184_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg935_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg36_out_to_MUX_Product106_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product106_3_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product106_3_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product107_3_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product107_3_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product107_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product107_3_impl_out,
                 X => Delay1No172_out_to_Product107_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product107_3_impl_parent_implementedSystem_port_1_cast);

SharedReg35_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg862_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg809_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg809_out;
SharedReg880_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg880_out;
SharedReg392_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg392_out;
SharedReg471_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg471_out;
SharedReg813_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg813_out;
SharedReg835_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg936_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg919_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg919_out;
SharedReg939_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg881_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg881_out;
   MUX_Product107_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg919_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg881_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg809_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg880_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg392_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg471_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg813_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg936_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product107_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product107_3_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product107_3_impl_0_out,
                 Y => Delay1No172_out);

SharedReg918_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg955_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg955_out;
SharedReg943_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg944_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg944_out;
SharedReg1002_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1002_out;
SharedReg183_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg183_out;
SharedReg982_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg982_out;
SharedReg1012_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1012_out;
SharedReg936_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg106_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg106_out;
SharedReg939_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg966_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg966_out;
   MUX_Product107_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg955_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg106_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg966_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg944_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1002_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg183_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg982_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1012_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg936_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product107_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product107_3_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product107_3_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product114_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_3_impl_out,
                 X => Delay1No174_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
Delay80No2_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast <= Delay80No2_out;
SharedReg864_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg864_out;
SharedReg140_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg512_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg512_out;
SharedReg470_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg470_out;
SharedReg829_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg398_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg398_out;
SharedReg581_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg581_out;
SharedReg937_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg674_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg674_out;
SharedReg939_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg665_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg665_out;
   MUX_Product114_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay80No2_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg674_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg665_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg864_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg140_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg512_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg470_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg398_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg581_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product114_3_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_3_impl_0_out,
                 Y => Delay1No174_out);

SharedReg941_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg941_out;
Delay81No9_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast <= Delay81No9_out;
SharedReg680_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg680_out;
SharedReg178_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg947_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg947_out;
SharedReg216_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg217_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg217_out;
SharedReg1014_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1014_out;
SharedReg951_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg937_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg147_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg147_out;
SharedReg939_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
SharedReg218_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg218_out;
   MUX_Product114_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay81No9_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg147_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg218_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg680_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg947_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg216_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg217_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1014_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product114_3_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_3_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product181_2_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product181_2_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product181_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product181_2_impl_out,
                 X => Delay1No176_out_to_Product181_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product181_2_impl_parent_implementedSystem_port_1_cast);

SharedReg682_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg682_out;
SharedReg53_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg309_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg309_out;
SharedReg849_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg849_out;
Delay1No218_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_5_cast <= Delay1No218_out;
SharedReg149_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg149_out;
SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg936_out;
SharedReg456_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg456_out;
SharedReg522_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg522_out;
SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg285_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg285_out;
SharedReg460_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg460_out;
SharedReg249_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg249_out;
   MUX_Product181_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg682_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg285_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg460_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg249_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg309_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay1No218_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg149_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg456_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg522_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product181_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product181_2_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_2_impl_0_out,
                 Y => Delay1No176_out);

SharedReg652_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg164_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg164_out;
SharedReg62_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg956_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg956_out;
SharedReg931_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg111_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg111_out;
SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg936_out;
SharedReg165_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg89_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg89_out;
SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg936_out;
SharedReg994_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg994_out;
SharedReg938_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg938_out;
SharedReg750_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg750_out;
   MUX_Product181_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg164_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg994_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg938_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg750_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg62_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg956_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg111_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg89_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg936_out_to_MUX_Product181_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product181_2_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_2_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product461_3_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product461_3_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product461_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product461_3_impl_out,
                 X => Delay1No178_out_to_Product461_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product461_3_impl_parent_implementedSystem_port_1_cast);

SharedReg68_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg870_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg870_out;
SharedReg182_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg182_out;
SharedReg881_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg881_out;
SharedReg932_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg932_out;
SharedReg588_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg588_out;
SharedReg212_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg212_out;
SharedReg566_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg566_out;
SharedReg542_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg542_out;
SharedReg937_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg863_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg863_out;
SharedReg664_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg664_out;
SharedReg884_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg884_out;
   MUX_Product461_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg870_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg863_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg664_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg884_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg182_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg881_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg932_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg588_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg212_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg566_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg542_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product461_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product461_3_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_3_impl_0_out,
                 Y => Delay1No178_out);

SharedReg181_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg968_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg968_out;
SharedReg718_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg718_out;
SharedReg957_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg957_out;
SharedReg932_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg932_out;
SharedReg981_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg981_out;
SharedReg141_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg141_out;
SharedReg992_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg992_out;
SharedReg70_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg70_out;
SharedReg937_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg937_out;
SharedReg975_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg975_out;
SharedReg723_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg723_out;
SharedReg966_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg966_out;
   MUX_Product461_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg968_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg975_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg723_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg966_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg718_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg957_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg932_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg981_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg141_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg992_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg70_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg937_out_to_MUX_Product461_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product461_3_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_3_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product68_3_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product68_3_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product68_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_3_impl_out,
                 X => Delay1No180_out_to_Product68_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product68_3_impl_parent_implementedSystem_port_1_cast);

SharedReg68_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg826_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg826_out;
SharedReg30_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg869_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg869_out;
SharedReg928_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg928_out;
SharedReg885_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg885_out;
SharedReg865_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg865_out;
SharedReg805_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg805_out;
SharedReg142_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg142_out;
Delay88No2_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_10_cast <= Delay88No2_out;
SharedReg881_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg881_out;
SharedReg833_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg833_out;
SharedReg67_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg67_out;
   MUX_Product68_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg826_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg881_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg833_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg67_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg30_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg869_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg928_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg885_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg865_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg805_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg142_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay88No2_out_to_MUX_Product68_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product68_3_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_3_impl_0_out,
                 Y => Delay1No180_out);

SharedReg215_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg955_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg955_out;
SharedReg139_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg957_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg957_out;
SharedReg945_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg945_out;
SharedReg981_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg981_out;
SharedReg934_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg934_out;
SharedReg961_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg961_out;
SharedReg213_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg213_out;
Delay100No_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_10_cast <= Delay100No_out;
SharedReg938_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg996_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg996_out;
SharedReg214_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg214_out;
   MUX_Product68_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg955_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg996_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg214_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg139_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg957_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg945_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg981_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg934_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg961_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg213_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay100No_out_to_MUX_Product68_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product68_3_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_3_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product911_3_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product911_3_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product911_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product911_3_impl_out,
                 X => Delay1No182_out_to_Product911_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product911_3_impl_parent_implementedSystem_port_1_cast);

SharedReg868_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg868_out;
SharedReg811_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg811_out;
SharedReg873_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg873_out;
SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg872_out;
SharedReg930_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg930_out;
SharedReg828_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg828_out;
SharedReg212_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg212_out;
SharedReg832_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg832_out;
SharedReg552_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg552_out;
SharedReg867_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg867_out;
SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg872_out;
SharedReg871_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg871_out;
SharedReg917_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg917_out;
   MUX_Product911_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg868_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg811_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg871_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg917_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg873_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg872_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg930_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg828_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg212_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg832_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg552_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg867_out_to_MUX_Product911_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product911_3_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_3_impl_0_out,
                 Y => Delay1No182_out);

SharedReg954_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg954_out;
SharedReg978_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg978_out;
SharedReg956_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg956_out;
SharedReg944_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg944_out;
SharedReg945_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg945_out;
SharedReg971_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg971_out;
SharedReg101_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg101_out;
SharedReg992_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg992_out;
SharedReg38_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg950_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg950_out;
SharedReg938_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg986_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg986_out;
SharedReg716_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg716_out;
   MUX_Product911_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg954_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg978_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg986_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg716_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg956_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg944_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg945_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg971_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg101_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg992_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg950_out_to_MUX_Product911_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product911_3_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_3_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product97_3_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product97_3_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product97_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product97_3_impl_out,
                 X => Delay1No184_out_to_Product97_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product97_3_impl_parent_implementedSystem_port_1_cast);

SharedReg35_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg34_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg34_out;
SharedReg66_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg179_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg179_out;
Delay14No10_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_5_cast <= Delay14No10_out;
Delay1No220_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_6_cast <= Delay1No220_out;
SharedReg859_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg859_out;
SharedReg788_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg788_out;
Delay50No_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_9_cast <= Delay50No_out;
SharedReg876_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg876_out;
SharedReg671_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg671_out;
SharedReg664_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg664_out;
   MUX_Product97_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg671_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg664_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg66_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg179_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay14No10_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay1No220_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg859_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg788_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay50No_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg876_out_to_MUX_Product97_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product97_3_impl_0_LUT_out,
                 oMux => MUX_Product97_3_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product97_3_impl_0_out,
                 Y => Delay1No184_out);

SharedReg104_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg100_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg143_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
SharedReg724_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg724_out;
SharedReg920_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg917_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg917_out;
SharedReg942_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg942_out;
SharedReg936_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg936_out;
SharedReg951_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg951_out;
SharedReg1004_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1004_out;
SharedReg943_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg943_out;
SharedReg931_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg931_out;
   MUX_Product97_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg943_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg931_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg143_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg724_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg917_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg942_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg936_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg951_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1004_out_to_MUX_Product97_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product97_3_impl_1_LUT_out,
                 oMux => MUX_Product97_3_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product97_3_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Subtract12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_0_impl_out,
                 X => Delay1No186_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg228_out;
SharedReg448_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg448_out;
Delay91No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast <= Delay91No_out;
SharedReg416_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg407_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg407_out;
SharedReg348_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg348_out;
SharedReg281_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg281_out;
SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg230_out;
SharedReg445_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg224_out;
SharedReg305_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg305_out;
SharedReg295_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg295_out;
   MUX_Subtract12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg224_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg305_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg295_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg448_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay91No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg407_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg348_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg281_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg230_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_0_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_0_out,
                 Y => Delay1No186_out);

SharedReg592_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg592_out;
SharedReg730_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg730_out;
SharedReg728_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg728_out;
SharedReg683_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg683_out;
SharedReg611_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg611_out;
Delay65No1_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast <= Delay65No1_out;
SharedReg739_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg739_out;
SharedReg702_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg702_out;
SharedReg733_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg733_out;
SharedReg732_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg732_out;
SharedReg590_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg590_out;
SharedReg734_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg734_out;
SharedReg589_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg589_out;
   MUX_Subtract12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg592_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg730_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg590_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg734_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg589_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg728_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg683_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg611_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay65No1_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg739_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg702_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg733_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg732_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_0_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Subtract12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_1_impl_out,
                 X => Delay1No188_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg534_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg377_out;
Delay73No_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast <= Delay73No_out;
SharedReg426_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg450_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg450_out;
SharedReg524_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg524_out;
SharedReg412_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg412_out;
SharedReg854_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg854_out;
SharedReg298_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg298_out;
SharedReg294_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg294_out;
SharedReg492_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg492_out;
SharedReg351_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg351_out;
   MUX_Subtract12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg294_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg492_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg351_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay73No_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg426_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg450_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg524_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg412_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg854_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg298_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_1_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_0_out,
                 Y => Delay1No188_out);

SharedReg638_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg638_out;
SharedReg596_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg653_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg653_out;
Delay63No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast <= Delay63No_out;
SharedReg659_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg659_out;
SharedReg612_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg612_out;
SharedReg606_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg606_out;
SharedReg683_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg683_out;
SharedReg620_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg620_out;
SharedReg594_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg594_out;
Delay40No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast <= Delay40No_out;
SharedReg739_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg739_out;
SharedReg684_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg684_out;
   MUX_Subtract12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg638_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay40No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg739_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg684_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg653_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay63No_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg659_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg612_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg606_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg683_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg620_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg594_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_1_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Subtract12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_2_impl_out,
                 X => Delay1No190_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg247_out;
Delay83No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast <= Delay83No5_out;
SharedReg583_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg583_out;
SharedReg280_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg280_out;
SharedReg804_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg804_out;
SharedReg286_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg354_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg354_out;
SharedReg512_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg512_out;
SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg374_out;
SharedReg432_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg432_out;
SharedReg473_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg473_out;
SharedReg838_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg838_out;
   MUX_Subtract12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg247_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg432_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg473_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg838_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay83No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg583_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg280_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg804_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg354_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg512_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_2_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_0_out,
                 Y => Delay1No190_out);

SharedReg618_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg618_out;
SharedReg704_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg704_out;
SharedReg699_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg699_out;
SharedReg757_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg757_out;
SharedReg715_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg715_out;
SharedReg638_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg638_out;
SharedReg747_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg747_out;
SharedReg706_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg706_out;
SharedReg742_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg742_out;
SharedReg710_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg710_out;
SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg623_out;
SharedReg721_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg721_out;
SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg623_out;
   MUX_Subtract12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg618_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg704_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg721_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg623_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg699_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg757_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg715_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg638_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg747_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg706_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg742_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg710_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_2_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Subtract1_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract1_3_impl_out,
                 X => Delay1No192_out_to_Subtract1_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Subtract1_3_impl_parent_implementedSystem_port_1_cast);

SharedReg571_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg357_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg327_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg327_out;
SharedReg570_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg834_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg834_out;
SharedReg478_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg478_out;
SharedReg383_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg383_out;
SharedReg292_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg292_out;
SharedReg792_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg792_out;
SharedReg565_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg565_out;
SharedReg839_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg839_out;
SharedReg805_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg805_out;
SharedReg866_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg866_out;
   MUX_Subtract1_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg839_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg805_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg866_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg327_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg834_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg478_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg383_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg292_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg792_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg565_out_to_MUX_Subtract1_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract1_3_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_3_impl_0_out,
                 Y => Delay1No192_out);

SharedReg743_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg743_out;
SharedReg662_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg662_out;
SharedReg714_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg714_out;
SharedReg719_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg719_out;
SharedReg756_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg756_out;
SharedReg664_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg664_out;
SharedReg619_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg619_out;
SharedReg621_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg621_out;
SharedReg720_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg720_out;
SharedReg616_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg616_out;
SharedReg712_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg712_out;
SharedReg671_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg671_out;
SharedReg748_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg748_out;
   MUX_Subtract1_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg743_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg662_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg712_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg671_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg748_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg714_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg719_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg756_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg664_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg619_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg621_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg720_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg616_out_to_MUX_Subtract1_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract1_3_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_3_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Add10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Add10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Add10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add10_3_impl_out,
                 X => Delay1No194_out_to_Add10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Add10_3_impl_parent_implementedSystem_port_1_cast);

Delay7No16_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_1_cast <= Delay7No16_out;
SharedReg868_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg868_out;
SharedReg874_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg874_out;
SharedReg875_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg875_out;
SharedReg860_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg860_out;
SharedReg857_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg857_out;
SharedReg867_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg867_out;
SharedReg873_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg873_out;
   MUX_Add10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No16_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg868_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg874_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg875_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg860_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg857_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg867_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg873_out_to_MUX_Add10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iSel => MUX_Add10_3_impl_0_LUT_out,
                 oMux => MUX_Add10_3_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_3_impl_0_out,
                 Y => Delay1No194_out);

SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg664_out;
SharedReg623_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg623_out;
SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg917_out;
SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg917_out;
SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg664_out;
SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg917_out;
SharedReg928_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg928_out;
   MUX_Add10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg623_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg664_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg917_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg928_out_to_MUX_Add10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iSel => MUX_Add10_3_impl_1_LUT_out,
                 oMux => MUX_Add10_3_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_3_impl_1_out,
                 Y => Delay1No195_out);
   Constant1_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

Delay1No196_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Divide_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_0_impl_out,
                 X => Delay1No196_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast);

SharedReg924_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg924_out;
SharedReg926_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg926_out;
SharedReg925_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg925_out;
Delay103No1_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast <= Delay103No1_out;
   MUX_Divide_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg924_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg925_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay103No1_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Divide_0_impl_0_LUT_out,
                 oMux => MUX_Divide_0_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_0_out,
                 Y => Delay1No196_out);

SharedReg727_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg727_out;
SharedReg652_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg652_out;
SharedReg711_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg711_out;
SharedReg716_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg716_out;
   MUX_Divide_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg727_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg652_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg711_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg716_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Divide_0_impl_1_LUT_out,
                 oMux => MUX_Divide_0_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product3_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product3_3_impl_out,
                 X => Delay1No198_out_to_Product3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
Delay1No224_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_2_cast <= Delay1No224_out;
Delay67No1_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_3_cast <= Delay67No1_out;
SharedReg928_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg928_out;
SharedReg872_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg872_out;
SharedReg880_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg880_out;
SharedReg667_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg667_out;
   MUX_Product3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No224_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay67No1_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg928_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg872_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg880_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg667_out_to_MUX_Product3_3_impl_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_Product3_3_impl_0_LUT_out,
                 oMux => MUX_Product3_3_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product3_3_impl_0_out,
                 Y => Delay1No198_out);

SharedReg102_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg102_out;
SharedReg220_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg220_out;
SharedReg941_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg941_out;
SharedReg959_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg959_out;
SharedReg948_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg948_out;
SharedReg1006_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1006_out;
SharedReg931_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg931_out;
   MUX_Product3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg102_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg220_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg941_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg959_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg948_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1006_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg931_out_to_MUX_Product3_3_impl_1_parent_implementedSystem_port_7_cast,
                 iSel => MUX_Product3_3_impl_1_LUT_out,
                 oMux => MUX_Product3_3_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product3_3_impl_1_out,
                 Y => Delay1No199_out);
   Constant_0_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);

   Delay16No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_0_out,
                 Y => Delay16No_out);

   Delay6No_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_1_out,
                 Y => Delay6No_out);

   Delay7No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_2_out,
                 Y => Delay7No_out);

   Delay19No_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_3_out,
                 Y => Delay19No_out);

   Delay103No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => Delay103No_out);

   Delay108No_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => Delay108No_out);

   Delay108No1_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => Delay108No1_out);

   Delay100No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay100No_out);

   Delay90No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay90No_out);

   Delay100No1_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => Delay100No1_out);

   Delay18No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => Delay18No2_out);

   Delay93No1_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => Delay93No1_out);

   Delay107No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => Delay107No_out);

   Delay111No_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => Delay111No_out);

   Delay100No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => Delay100No2_out);

   Delay96No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => Delay96No2_out);

   Delay3No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_0_out,
                 Y => Delay3No2_out);

   Delay6No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_1_out,
                 Y => Delay6No4_out);

   Delay4No7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_2_out,
                 Y => Delay4No7_out);

   Delay7No7_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_3_out,
                 Y => Delay7No7_out);

   Delay87No_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => Delay87No_out);

   Delay94No1_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay94No1_out);

   Delay108No2_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay108No2_out);

   Delay107No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => Delay107No1_out);

   Delay93No2_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => Delay93No2_out);

   Delay80No1_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => Delay80No1_out);

   Delay93No3_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => Delay93No3_out);

   Delay97No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => Delay97No_out);

   Delay94No3_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => Delay94No3_out);

   Delay93No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => Delay93No4_out);

   Delay90No1_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => Delay90No1_out);

   Delay87No3_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => Delay87No3_out);

   Delay3No10_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_0_out,
                 Y => Delay3No10_out);

   Delay6No9_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_1_out,
                 Y => Delay6No9_out);

   Delay4No9_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_2_out,
                 Y => Delay4No9_out);

   Delay7No16_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_3_out,
                 Y => Delay7No16_out);

   Delay12No12_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_0_out,
                 Y => Delay12No12_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_1_out,
                 Y => Delay1No215_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_2_out,
                 Y => Delay1No216_out);

   Delay14No10_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_3_out,
                 Y => Delay14No10_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_0_out,
                 Y => Delay1No217_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_1_out,
                 Y => Delay1No218_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_2_out,
                 Y => Delay1No219_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_3_out,
                 Y => Delay1No220_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_0_out,
                 Y => Delay1No221_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_1_out,
                 Y => Delay1No222_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_2_out,
                 Y => Delay1No223_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_3_out,
                 Y => Delay1No224_out);

   Delay65No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => Delay65No1_out);

   Delay12No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => Delay12No15_out);

   Delay63No_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => Delay63No_out);

   Delay59No_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => Delay59No_out);

   Delay84No1_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => Delay84No1_out);

   Delay40No_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => Delay40No_out);

   Delay96No3_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => Delay96No3_out);

   Delay96No4_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => Delay96No4_out);

   Delay79No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => Delay79No_out);

   Delay80No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => Delay80No2_out);

   Delay58No1_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => Delay58No1_out);

   Delay87No5_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => Delay87No5_out);

   Delay73No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => Delay73No_out);

   Delay77No2_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => Delay77No2_out);

   Delay75No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => Delay75No1_out);

   Delay83No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => Delay83No4_out);

   Delay91No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => Delay91No_out);

   Delay94No4_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => Delay94No4_out);

   Delay98No_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => Delay98No_out);

   Delay94No5_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => Delay94No5_out);

   Delay97No1_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => Delay97No1_out);

   Delay87No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => Delay87No6_out);

   Delay76No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay76No2_out);

   Delay93No5_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => Delay93No5_out);

   Delay93No6_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => Delay93No6_out);

   Delay98No1_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => Delay98No1_out);

   Delay89No1_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => Delay89No1_out);

   Delay85No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => Delay85No2_out);

   Delay94No6_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => Delay94No6_out);

   Delay79No4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => Delay79No4_out);

   Delay83No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => Delay83No5_out);

   Delay78No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => Delay78No1_out);

   Delay95No_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => Delay95No_out);

   Delay99No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => Delay99No1_out);

   Delay87No7_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => Delay87No7_out);

   Delay90No2_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => Delay90No2_out);

   Delay85No3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => Delay85No3_out);

   Delay89No2_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => Delay89No2_out);

   Delay68No3_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => Delay68No3_out);

   Delay101No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => Delay101No_out);

   Delay82No6_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => Delay82No6_out);

   Delay92No_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => Delay92No_out);

   Delay88No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => Delay88No2_out);

   Delay90No3_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => Delay90No3_out);

   Delay82No7_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => Delay82No7_out);

   Delay84No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => Delay84No4_out);

   Delay79No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => Delay79No5_out);

   Delay85No4_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay85No4_out);

   Delay68No4_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => Delay68No4_out);

   Delay85No5_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => Delay85No5_out);

   Delay96No6_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => Delay96No6_out);

   Delay56No3_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay56No3_out);

   Delay48No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => Delay48No_out);

   Delay90No4_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => Delay90No4_out);

   Delay79No7_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => Delay79No7_out);

   Delay87No8_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => Delay87No8_out);

   Delay13No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => Delay13No41_out);

   Delay73No2_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => Delay73No2_out);

   Delay79No8_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => Delay79No8_out);

   Delay103No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => Delay103No1_out);

   Delay54No_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => Delay54No_out);

   Delay50No_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => Delay50No_out);

   Delay64No4_instance: Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=51 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => Delay64No4_out);

   Delay67No1_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => Delay67No1_out);

   Delay71No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => Delay71No6_out);

   Delay97No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => Delay97No2_out);

   Delay97No3_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => Delay97No3_out);

   Delay98No2_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => Delay98No2_out);

   Delay86No6_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => Delay86No6_out);

   Delay96No7_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => Delay96No7_out);

   Delay81No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => Delay81No8_out);

   Delay80No9_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => Delay80No9_out);

   Delay81No9_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => Delay81No9_out);

   Delay100No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => Delay100No4_out);

   MUX_Add121_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add121_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add121_3_impl_0_LUT_out);

   MUX_Add121_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add121_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add121_3_impl_1_LUT_out);

   MUX_Add22_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add22_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add22_3_impl_0_LUT_out);

   MUX_Add22_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add22_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add22_3_impl_1_LUT_out);

   MUX_Product97_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product97_3_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product97_3_impl_0_LUT_out);

   MUX_Product97_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product97_3_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product97_3_impl_1_LUT_out);

   MUX_Add10_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add10_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add10_3_impl_0_LUT_out);

   MUX_Add10_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add10_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add10_3_impl_1_LUT_out);

   MUX_Divide_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Divide_0_impl_0_LUT_out);

   MUX_Divide_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Divide_0_impl_1_LUT_out);

   MUX_Product3_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product3_3_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product3_3_impl_0_LUT_out);

   MUX_Product3_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product3_3_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product3_3_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=86 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_1_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_2_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_3_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_0_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_1_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_2_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_3_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_0_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_1_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_2_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_3_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_0_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_1_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_2_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_3_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_0_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_1_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_2_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=59 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_3_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_0_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_1_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_2_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_3_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_0_impl_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_1_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_2_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_3_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_0_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_1_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_2_impl_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_3_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_0_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=59 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_1_impl_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_2_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_3_impl_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_0_impl_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_1_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_2_impl_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_3_impl_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_0_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_1_impl_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_2_impl_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_3_impl_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_0_impl_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_1_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_2_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_3_impl_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_0_impl_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_1_impl_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_2_impl_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_3_impl_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_0_impl_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_1_impl_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_2_impl_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_3_impl_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_1_impl_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_3_impl_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_1_impl_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_3_impl_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_1_impl_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_3_impl_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_1_impl_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_3_impl_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_0_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_1_impl_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_2_impl_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_3_impl_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_1_impl_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_2_impl_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_3_impl_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_1_impl_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_1_impl_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_2_impl_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_3_impl_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_0_impl_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_1_impl_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add17_3_impl_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add22_3_impl_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_1_impl_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_2_impl_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_2_impl_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_3_impl_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product103_2_impl_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product103_3_impl_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product106_3_impl_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product107_3_impl_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_3_impl_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product181_2_impl_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product461_3_impl_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg857_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_3_impl_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product911_3_impl_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product97_3_impl_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_0_impl_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_1_impl_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_2_impl_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract1_3_impl_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add10_3_impl_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg918_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_0_impl_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product3_3_impl_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg934_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg938_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg965_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg967_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg971_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg983_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg984_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg985_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg997_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1000_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1003_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1006_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1010_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);
end architecture;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity implementedSystem_toplevel_wrapper is
  port (
    clk, rst : in std_logic;
    shared_input : in std_logic_vector(31 downto 0);
    ldiff_uu_del_1_0_enable : in std_logic;
    ldiff_uu_del_1_1_enable : in std_logic;
    ldiff_uu_del_1_2_enable : in std_logic;
    ldiff_uu_del_1_3_enable : in std_logic;
    ldiff_uv_del_1_0_enable : in std_logic;
    ldiff_uv_del_1_1_enable : in std_logic;
    ldiff_uv_del_1_2_enable : in std_logic;
    ldiff_uv_del_1_3_enable : in std_logic;
    ldiff_uw_del_1_0_enable : in std_logic;
    ldiff_uw_del_1_1_enable : in std_logic;
    ldiff_uw_del_1_2_enable : in std_logic;
    ldiff_uw_del_1_3_enable : in std_logic;
    ldiff_vu_del_1_0_enable : in std_logic;
    ldiff_vu_del_1_1_enable : in std_logic;
    ldiff_vu_del_1_2_enable : in std_logic;
    ldiff_vu_del_1_3_enable : in std_logic;
    ldiff_vv_del_1_0_enable : in std_logic;
    ldiff_vv_del_1_1_enable : in std_logic;
    ldiff_vv_del_1_2_enable : in std_logic;
    ldiff_vv_del_1_3_enable : in std_logic;
    ldiff_vw_del_1_0_enable : in std_logic;
    ldiff_vw_del_1_1_enable : in std_logic;
    ldiff_vw_del_1_2_enable : in std_logic;
    ldiff_vw_del_1_3_enable : in std_logic;
    ldiff_wu_del_1_0_enable : in std_logic;
    ldiff_wu_del_1_1_enable : in std_logic;
    ldiff_wu_del_1_2_enable : in std_logic;
    ldiff_wu_del_1_3_enable : in std_logic;
    ldiff_wv_del_1_0_enable : in std_logic;
    ldiff_wv_del_1_1_enable : in std_logic;
    ldiff_wv_del_1_2_enable : in std_logic;
    ldiff_wv_del_1_3_enable : in std_logic;
    ldiff_ww_del_1_0_enable : in std_logic;
    ldiff_ww_del_1_1_enable : in std_logic;
    ldiff_ww_del_1_2_enable : in std_logic;
    ldiff_ww_del_1_3_enable : in std_logic;
    r_u_0_enable : in std_logic;
    r_u_1_enable : in std_logic;
    r_u_2_enable : in std_logic;
    r_u_3_enable : in std_logic;
    r_v_0_enable : in std_logic;
    r_v_1_enable : in std_logic;
    r_v_2_enable : in std_logic;
    r_v_3_enable : in std_logic;
    r_w_0_enable : in std_logic;
    r_w_1_enable : in std_logic;
    r_w_2_enable : in std_logic;
    r_w_3_enable : in std_logic;
    output_select : in std_logic_vector(5 downto 0);
    shared_output : out std_logic_vector(31 downto 0)
  );
end entity;

architecture implementedSystem_toplevel_wrapper of implementedSystem_toplevel_wrapper is
  signal ldiff_uu_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uu_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uu_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uu_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uv_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uv_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uv_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uv_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uw_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uw_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uw_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_uw_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vu_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vu_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vu_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vu_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vv_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vv_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vv_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vv_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vw_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vw_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vw_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_vw_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wu_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wu_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wu_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wu_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wv_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wv_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wv_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_wv_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_ww_del_1_0_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_ww_del_1_1_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_ww_del_1_2_DUT_in : std_logic_vector(31 downto 0);
  signal ldiff_ww_del_1_3_DUT_in : std_logic_vector(31 downto 0);
  signal r_u_0_DUT_in : std_logic_vector(31 downto 0);
  signal r_u_1_DUT_in : std_logic_vector(31 downto 0);
  signal r_u_2_DUT_in : std_logic_vector(31 downto 0);
  signal r_u_3_DUT_in : std_logic_vector(31 downto 0);
  signal r_v_0_DUT_in : std_logic_vector(31 downto 0);
  signal r_v_1_DUT_in : std_logic_vector(31 downto 0);
  signal r_v_2_DUT_in : std_logic_vector(31 downto 0);
  signal r_v_3_DUT_in : std_logic_vector(31 downto 0);
  signal r_w_0_DUT_in : std_logic_vector(31 downto 0);
  signal r_w_1_DUT_in : std_logic_vector(31 downto 0);
  signal r_w_2_DUT_in : std_logic_vector(31 downto 0);
  signal r_w_3_DUT_in : std_logic_vector(31 downto 0);
  signal inv_11_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_11_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_11_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_11_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_12_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_12_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_12_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_12_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_13_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_13_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_13_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_13_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_21_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_21_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_21_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_21_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_22_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_22_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_22_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_22_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_23_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_23_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_23_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_23_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_31_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_31_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_31_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_31_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_32_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_32_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_32_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_32_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_33_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_33_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_33_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_33_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_41_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_41_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_41_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_41_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_42_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_42_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_42_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_42_3_DUT_out : std_logic_vector(31 downto 0);
  signal inv_43_0_DUT_out : std_logic_vector(31 downto 0);
  signal inv_43_1_DUT_out : std_logic_vector(31 downto 0);
  signal inv_43_2_DUT_out : std_logic_vector(31 downto 0);
  signal inv_43_3_DUT_out : std_logic_vector(31 downto 0);
  type output_mux_input_t is array (0 to 47) of std_logic_vector(31 downto 0);
  signal output_mux_input : output_mux_input_t;

  begin
    DUT : entity work.implementedSystem_toplevel
      port map (
        clk => clk,
        rst => rst,
        ldiff_uu_del_1_0 => ldiff_uu_del_1_0_DUT_in,
        ldiff_uu_del_1_1 => ldiff_uu_del_1_1_DUT_in,
        ldiff_uu_del_1_2 => ldiff_uu_del_1_2_DUT_in,
        ldiff_uu_del_1_3 => ldiff_uu_del_1_3_DUT_in,
        ldiff_uv_del_1_0 => ldiff_uv_del_1_0_DUT_in,
        ldiff_uv_del_1_1 => ldiff_uv_del_1_1_DUT_in,
        ldiff_uv_del_1_2 => ldiff_uv_del_1_2_DUT_in,
        ldiff_uv_del_1_3 => ldiff_uv_del_1_3_DUT_in,
        ldiff_uw_del_1_0 => ldiff_uw_del_1_0_DUT_in,
        ldiff_uw_del_1_1 => ldiff_uw_del_1_1_DUT_in,
        ldiff_uw_del_1_2 => ldiff_uw_del_1_2_DUT_in,
        ldiff_uw_del_1_3 => ldiff_uw_del_1_3_DUT_in,
        ldiff_vu_del_1_0 => ldiff_vu_del_1_0_DUT_in,
        ldiff_vu_del_1_1 => ldiff_vu_del_1_1_DUT_in,
        ldiff_vu_del_1_2 => ldiff_vu_del_1_2_DUT_in,
        ldiff_vu_del_1_3 => ldiff_vu_del_1_3_DUT_in,
        ldiff_vv_del_1_0 => ldiff_vv_del_1_0_DUT_in,
        ldiff_vv_del_1_1 => ldiff_vv_del_1_1_DUT_in,
        ldiff_vv_del_1_2 => ldiff_vv_del_1_2_DUT_in,
        ldiff_vv_del_1_3 => ldiff_vv_del_1_3_DUT_in,
        ldiff_vw_del_1_0 => ldiff_vw_del_1_0_DUT_in,
        ldiff_vw_del_1_1 => ldiff_vw_del_1_1_DUT_in,
        ldiff_vw_del_1_2 => ldiff_vw_del_1_2_DUT_in,
        ldiff_vw_del_1_3 => ldiff_vw_del_1_3_DUT_in,
        ldiff_wu_del_1_0 => ldiff_wu_del_1_0_DUT_in,
        ldiff_wu_del_1_1 => ldiff_wu_del_1_1_DUT_in,
        ldiff_wu_del_1_2 => ldiff_wu_del_1_2_DUT_in,
        ldiff_wu_del_1_3 => ldiff_wu_del_1_3_DUT_in,
        ldiff_wv_del_1_0 => ldiff_wv_del_1_0_DUT_in,
        ldiff_wv_del_1_1 => ldiff_wv_del_1_1_DUT_in,
        ldiff_wv_del_1_2 => ldiff_wv_del_1_2_DUT_in,
        ldiff_wv_del_1_3 => ldiff_wv_del_1_3_DUT_in,
        ldiff_ww_del_1_0 => ldiff_ww_del_1_0_DUT_in,
        ldiff_ww_del_1_1 => ldiff_ww_del_1_1_DUT_in,
        ldiff_ww_del_1_2 => ldiff_ww_del_1_2_DUT_in,
        ldiff_ww_del_1_3 => ldiff_ww_del_1_3_DUT_in,
        r_u_0 => r_u_0_DUT_in,
        r_u_1 => r_u_1_DUT_in,
        r_u_2 => r_u_2_DUT_in,
        r_u_3 => r_u_3_DUT_in,
        r_v_0 => r_v_0_DUT_in,
        r_v_1 => r_v_1_DUT_in,
        r_v_2 => r_v_2_DUT_in,
        r_v_3 => r_v_3_DUT_in,
        r_w_0 => r_w_0_DUT_in,
        r_w_1 => r_w_1_DUT_in,
        r_w_2 => r_w_2_DUT_in,
        r_w_3 => r_w_3_DUT_in,
        inv_11_0 => inv_11_0_DUT_out,
        inv_11_1 => inv_11_1_DUT_out,
        inv_11_2 => inv_11_2_DUT_out,
        inv_11_3 => inv_11_3_DUT_out,
        inv_12_0 => inv_12_0_DUT_out,
        inv_12_1 => inv_12_1_DUT_out,
        inv_12_2 => inv_12_2_DUT_out,
        inv_12_3 => inv_12_3_DUT_out,
        inv_13_0 => inv_13_0_DUT_out,
        inv_13_1 => inv_13_1_DUT_out,
        inv_13_2 => inv_13_2_DUT_out,
        inv_13_3 => inv_13_3_DUT_out,
        inv_21_0 => inv_21_0_DUT_out,
        inv_21_1 => inv_21_1_DUT_out,
        inv_21_2 => inv_21_2_DUT_out,
        inv_21_3 => inv_21_3_DUT_out,
        inv_22_0 => inv_22_0_DUT_out,
        inv_22_1 => inv_22_1_DUT_out,
        inv_22_2 => inv_22_2_DUT_out,
        inv_22_3 => inv_22_3_DUT_out,
        inv_23_0 => inv_23_0_DUT_out,
        inv_23_1 => inv_23_1_DUT_out,
        inv_23_2 => inv_23_2_DUT_out,
        inv_23_3 => inv_23_3_DUT_out,
        inv_31_0 => inv_31_0_DUT_out,
        inv_31_1 => inv_31_1_DUT_out,
        inv_31_2 => inv_31_2_DUT_out,
        inv_31_3 => inv_31_3_DUT_out,
        inv_32_0 => inv_32_0_DUT_out,
        inv_32_1 => inv_32_1_DUT_out,
        inv_32_2 => inv_32_2_DUT_out,
        inv_32_3 => inv_32_3_DUT_out,
        inv_33_0 => inv_33_0_DUT_out,
        inv_33_1 => inv_33_1_DUT_out,
        inv_33_2 => inv_33_2_DUT_out,
        inv_33_3 => inv_33_3_DUT_out,
        inv_41_0 => inv_41_0_DUT_out,
        inv_41_1 => inv_41_1_DUT_out,
        inv_41_2 => inv_41_2_DUT_out,
        inv_41_3 => inv_41_3_DUT_out,
        inv_42_0 => inv_42_0_DUT_out,
        inv_42_1 => inv_42_1_DUT_out,
        inv_42_2 => inv_42_2_DUT_out,
        inv_42_3 => inv_42_3_DUT_out,
        inv_43_0 => inv_43_0_DUT_out,
        inv_43_1 => inv_43_1_DUT_out,
        inv_43_2 => inv_43_2_DUT_out,
        inv_43_3 => inv_43_3_DUT_out
       );
    process(clk)
      begin
        if (rising_edge(clk)) then
          if (ldiff_uu_del_1_0_enable = '1') then
            ldiff_uu_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uu_del_1_0
          if (ldiff_uu_del_1_1_enable = '1') then
            ldiff_uu_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uu_del_1_1
          if (ldiff_uu_del_1_2_enable = '1') then
            ldiff_uu_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uu_del_1_2
          if (ldiff_uu_del_1_3_enable = '1') then
            ldiff_uu_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uu_del_1_3
          if (ldiff_uv_del_1_0_enable = '1') then
            ldiff_uv_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uv_del_1_0
          if (ldiff_uv_del_1_1_enable = '1') then
            ldiff_uv_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uv_del_1_1
          if (ldiff_uv_del_1_2_enable = '1') then
            ldiff_uv_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uv_del_1_2
          if (ldiff_uv_del_1_3_enable = '1') then
            ldiff_uv_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uv_del_1_3
          if (ldiff_uw_del_1_0_enable = '1') then
            ldiff_uw_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uw_del_1_0
          if (ldiff_uw_del_1_1_enable = '1') then
            ldiff_uw_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uw_del_1_1
          if (ldiff_uw_del_1_2_enable = '1') then
            ldiff_uw_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uw_del_1_2
          if (ldiff_uw_del_1_3_enable = '1') then
            ldiff_uw_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_uw_del_1_3
          if (ldiff_vu_del_1_0_enable = '1') then
            ldiff_vu_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vu_del_1_0
          if (ldiff_vu_del_1_1_enable = '1') then
            ldiff_vu_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vu_del_1_1
          if (ldiff_vu_del_1_2_enable = '1') then
            ldiff_vu_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vu_del_1_2
          if (ldiff_vu_del_1_3_enable = '1') then
            ldiff_vu_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vu_del_1_3
          if (ldiff_vv_del_1_0_enable = '1') then
            ldiff_vv_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vv_del_1_0
          if (ldiff_vv_del_1_1_enable = '1') then
            ldiff_vv_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vv_del_1_1
          if (ldiff_vv_del_1_2_enable = '1') then
            ldiff_vv_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vv_del_1_2
          if (ldiff_vv_del_1_3_enable = '1') then
            ldiff_vv_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vv_del_1_3
          if (ldiff_vw_del_1_0_enable = '1') then
            ldiff_vw_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vw_del_1_0
          if (ldiff_vw_del_1_1_enable = '1') then
            ldiff_vw_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vw_del_1_1
          if (ldiff_vw_del_1_2_enable = '1') then
            ldiff_vw_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vw_del_1_2
          if (ldiff_vw_del_1_3_enable = '1') then
            ldiff_vw_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_vw_del_1_3
          if (ldiff_wu_del_1_0_enable = '1') then
            ldiff_wu_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wu_del_1_0
          if (ldiff_wu_del_1_1_enable = '1') then
            ldiff_wu_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wu_del_1_1
          if (ldiff_wu_del_1_2_enable = '1') then
            ldiff_wu_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wu_del_1_2
          if (ldiff_wu_del_1_3_enable = '1') then
            ldiff_wu_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wu_del_1_3
          if (ldiff_wv_del_1_0_enable = '1') then
            ldiff_wv_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wv_del_1_0
          if (ldiff_wv_del_1_1_enable = '1') then
            ldiff_wv_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wv_del_1_1
          if (ldiff_wv_del_1_2_enable = '1') then
            ldiff_wv_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wv_del_1_2
          if (ldiff_wv_del_1_3_enable = '1') then
            ldiff_wv_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_wv_del_1_3
          if (ldiff_ww_del_1_0_enable = '1') then
            ldiff_ww_del_1_0_DUT_in <= shared_input;
          end if; -- enable for input ldiff_ww_del_1_0
          if (ldiff_ww_del_1_1_enable = '1') then
            ldiff_ww_del_1_1_DUT_in <= shared_input;
          end if; -- enable for input ldiff_ww_del_1_1
          if (ldiff_ww_del_1_2_enable = '1') then
            ldiff_ww_del_1_2_DUT_in <= shared_input;
          end if; -- enable for input ldiff_ww_del_1_2
          if (ldiff_ww_del_1_3_enable = '1') then
            ldiff_ww_del_1_3_DUT_in <= shared_input;
          end if; -- enable for input ldiff_ww_del_1_3
          if (r_u_0_enable = '1') then
            r_u_0_DUT_in <= shared_input;
          end if; -- enable for input r_u_0
          if (r_u_1_enable = '1') then
            r_u_1_DUT_in <= shared_input;
          end if; -- enable for input r_u_1
          if (r_u_2_enable = '1') then
            r_u_2_DUT_in <= shared_input;
          end if; -- enable for input r_u_2
          if (r_u_3_enable = '1') then
            r_u_3_DUT_in <= shared_input;
          end if; -- enable for input r_u_3
          if (r_v_0_enable = '1') then
            r_v_0_DUT_in <= shared_input;
          end if; -- enable for input r_v_0
          if (r_v_1_enable = '1') then
            r_v_1_DUT_in <= shared_input;
          end if; -- enable for input r_v_1
          if (r_v_2_enable = '1') then
            r_v_2_DUT_in <= shared_input;
          end if; -- enable for input r_v_2
          if (r_v_3_enable = '1') then
            r_v_3_DUT_in <= shared_input;
          end if; -- enable for input r_v_3
          if (r_w_0_enable = '1') then
            r_w_0_DUT_in <= shared_input;
          end if; -- enable for input r_w_0
          if (r_w_1_enable = '1') then
            r_w_1_DUT_in <= shared_input;
          end if; -- enable for input r_w_1
          if (r_w_2_enable = '1') then
            r_w_2_DUT_in <= shared_input;
          end if; -- enable for input r_w_2
          if (r_w_3_enable = '1') then
            r_w_3_DUT_in <= shared_input;
          end if; -- enable for input r_w_3
        end if; -- clk
      end process;
    output_mux_input(0) <= inv_11_0_DUT_out;
    output_mux_input(1) <= inv_11_1_DUT_out;
    output_mux_input(2) <= inv_11_2_DUT_out;
    output_mux_input(3) <= inv_11_3_DUT_out;
    output_mux_input(4) <= inv_12_0_DUT_out;
    output_mux_input(5) <= inv_12_1_DUT_out;
    output_mux_input(6) <= inv_12_2_DUT_out;
    output_mux_input(7) <= inv_12_3_DUT_out;
    output_mux_input(8) <= inv_13_0_DUT_out;
    output_mux_input(9) <= inv_13_1_DUT_out;
    output_mux_input(10) <= inv_13_2_DUT_out;
    output_mux_input(11) <= inv_13_3_DUT_out;
    output_mux_input(12) <= inv_21_0_DUT_out;
    output_mux_input(13) <= inv_21_1_DUT_out;
    output_mux_input(14) <= inv_21_2_DUT_out;
    output_mux_input(15) <= inv_21_3_DUT_out;
    output_mux_input(16) <= inv_22_0_DUT_out;
    output_mux_input(17) <= inv_22_1_DUT_out;
    output_mux_input(18) <= inv_22_2_DUT_out;
    output_mux_input(19) <= inv_22_3_DUT_out;
    output_mux_input(20) <= inv_23_0_DUT_out;
    output_mux_input(21) <= inv_23_1_DUT_out;
    output_mux_input(22) <= inv_23_2_DUT_out;
    output_mux_input(23) <= inv_23_3_DUT_out;
    output_mux_input(24) <= inv_31_0_DUT_out;
    output_mux_input(25) <= inv_31_1_DUT_out;
    output_mux_input(26) <= inv_31_2_DUT_out;
    output_mux_input(27) <= inv_31_3_DUT_out;
    output_mux_input(28) <= inv_32_0_DUT_out;
    output_mux_input(29) <= inv_32_1_DUT_out;
    output_mux_input(30) <= inv_32_2_DUT_out;
    output_mux_input(31) <= inv_32_3_DUT_out;
    output_mux_input(32) <= inv_33_0_DUT_out;
    output_mux_input(33) <= inv_33_1_DUT_out;
    output_mux_input(34) <= inv_33_2_DUT_out;
    output_mux_input(35) <= inv_33_3_DUT_out;
    output_mux_input(36) <= inv_41_0_DUT_out;
    output_mux_input(37) <= inv_41_1_DUT_out;
    output_mux_input(38) <= inv_41_2_DUT_out;
    output_mux_input(39) <= inv_41_3_DUT_out;
    output_mux_input(40) <= inv_42_0_DUT_out;
    output_mux_input(41) <= inv_42_1_DUT_out;
    output_mux_input(42) <= inv_42_2_DUT_out;
    output_mux_input(43) <= inv_42_3_DUT_out;
    output_mux_input(44) <= inv_43_0_DUT_out;
    output_mux_input(45) <= inv_43_1_DUT_out;
    output_mux_input(46) <= inv_43_2_DUT_out;
    output_mux_input(47) <= inv_43_3_DUT_out;
    shared_output <= output_mux_input(to_integer(unsigned(output_select)));
    
end architecture;
