--------------------------------------------------------------------------------
--                         ModuloCounter_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_28_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of ModuloCounter_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(4 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 27 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_9_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2436208_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2436210)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2436208_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2436208_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2436213
--                  (IntAdderAlternative_27_f250_uid2436217)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2436213 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2436213 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2436220
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2436220 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2436220 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2436223
--                   (IntAdderClassical_34_f250_uid2436225)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2436223 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2436223 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2436208
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2436208 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2436208 is
   component FPAdd_8_23_uid2436208_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2436213 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2436220 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2436223 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2436208_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2436213  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2436220  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2436223  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2436208 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2436208  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_28_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_28_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_28_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
         iS_23 when "10111",
         iS_24 when "11000",
         iS_25 when "11001",
         iS_26 when "11010",
         iS_27 when "11011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2437397
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2437397 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2437397 is
signal XX_m2437398 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2437398 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2437398 <= X ;
   YY_m2437398 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2437401
--                   (IntAdderClassical_33_f500_uid2437403)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2437401 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2437401 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2437397 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2437401 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2437397  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2437401  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2437836_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2437838)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2437836_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2437836_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2437841
--                  (IntAdderAlternative_27_f250_uid2437845)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2437841 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2437841 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2437848
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2437848 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2437848 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2437851
--                   (IntAdderClassical_34_f250_uid2437853)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2437851 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2437851 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2437836
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2437836 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2437836 is
   component FPAdd_8_23_uid2437836_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2437841 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2437848 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2437851 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2437836_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2437841  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2437848  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2437851  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2437836 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2437836  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_20_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_20_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_20_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0010" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0011" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0100" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0101" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0110" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0111" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "1000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0001" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0010" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0011" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0100" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0101" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0110" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0111" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "1000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0001" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0110" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0111" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "1000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0001" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0010" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0011" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0100" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0101" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0001" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0010" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0011" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0100" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0101" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0011" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0100" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0101" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0110" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0111" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "1000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0001" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0010" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0101" when "00001",
      "0000" when "00010",
      "0000" when "00011",
      "0110" when "00100",
      "0000" when "00101",
      "0000" when "00110",
      "0111" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "1000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0001" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0010" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0011" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0100" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0101" when "00001",
      "0000" when "00010",
      "0000" when "00011",
      "0110" when "00100",
      "0000" when "00101",
      "0000" when "00110",
      "0111" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "1000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0001" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0010" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0011" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0100" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0001" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0010" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0011" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0100" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0101" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0110" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0111" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "1000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "1000" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0001" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0010" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0011" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0100" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0101" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0110" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0111" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0101" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0001" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0010" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0011" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0100" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0101" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0001" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0010" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0011" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0100" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0011" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0100" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0101" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0110" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0111" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "1000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0001" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0010" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0010" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0011" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0100" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0101" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0110" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0111" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "1000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0001" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0010" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0011" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0100" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0101" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0110" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0111" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "1000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0001" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0100" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0101" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0001" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0110" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0111" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "1000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0010" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0011" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0110" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0111" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "1000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0001" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0010" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0011" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0100" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0101" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0101" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0001" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0010" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0011" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0100" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0011" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0100" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0101" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0110" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0111" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "1000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0001" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0010" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0011" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0100" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0101" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0110" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0111" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "1000" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0001" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0010" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0101" when "00001",
      "0000" when "00010",
      "0000" when "00011",
      "0110" when "00100",
      "0000" when "00101",
      "0000" when "00110",
      "0111" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "1000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0001" when "10001",
      "0000" when "10010",
      "0000" when "10011",
      "0010" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0011" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0100" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0001" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0010" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0011" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0100" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0101" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0110" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0111" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "1000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0001" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0010" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0011" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0100" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0101" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0110" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0111" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "1000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0101" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0001" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0010" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0011" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0100" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0101" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0110" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0111" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0000" when "01001",
      "1000" when "01010",
      "0000" when "01011",
      "0000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0001" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "0010" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0011" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0100" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0010" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0011" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0100" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0101" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0110" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0111" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "1000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0001" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0010" when "00000",
      "0000" when "00001",
      "0000" when "00010",
      "0011" when "00011",
      "0000" when "00100",
      "0000" when "00101",
      "0100" when "00110",
      "0000" when "00111",
      "0000" when "01000",
      "0101" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "0110" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0111" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0000" when "10010",
      "1000" when "10011",
      "0000" when "10100",
      "0000" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0000" when "11000",
      "0001" when "11001",
      "0000" when "11010",
      "0000" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "0000" when "00000",
      "0000" when "00001",
      "0101" when "00010",
      "0000" when "00011",
      "0000" when "00100",
      "0110" when "00101",
      "0000" when "00110",
      "0000" when "00111",
      "0111" when "01000",
      "0000" when "01001",
      "0000" when "01010",
      "0000" when "01011",
      "1000" when "01100",
      "0000" when "01101",
      "0000" when "01110",
      "0000" when "01111",
      "0000" when "10000",
      "0000" when "10001",
      "0001" when "10010",
      "0000" when "10011",
      "0000" when "10100",
      "0010" when "10101",
      "0000" when "10110",
      "0000" when "10111",
      "0011" when "11000",
      "0000" when "11001",
      "0000" when "11010",
      "0100" when "11011",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "01011" when "00000",
      "01101" when "00001",
      "00000" when "00010",
      "00010" when "00011",
      "10000" when "00100",
      "00000" when "00101",
      "10011" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "10001" when "01001",
      "10010" when "01010",
      "00000" when "01011",
      "01110" when "01100",
      "01001" when "01101",
      "00000" when "01110",
      "00111" when "01111",
      "00110" when "10000",
      "00000" when "10001",
      "01111" when "10010",
      "01000" when "10011",
      "00001" when "10100",
      "00101" when "10101",
      "00011" when "10110",
      "01100" when "10111",
      "00000" when "11000",
      "01010" when "11001",
      "00100" when "11010",
      "00000" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5 is
signal t_in : std_logic_vector(4 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   with t_in select t_out <= 
      "00101" when "00000",
      "00110" when "00001",
      "00000" when "00010",
      "10011" when "00011",
      "00010" when "00100",
      "00000" when "00101",
      "00100" when "00110",
      "10010" when "00111",
      "00000" when "01000",
      "00011" when "01001",
      "00001" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "10000" when "01101",
      "00000" when "01110",
      "01111" when "01111",
      "01100" when "10000",
      "00000" when "10001",
      "01000" when "10010",
      "10001" when "10011",
      "01101" when "10100",
      "01110" when "10101",
      "01001" when "10110",
      "00111" when "10111",
      "00000" when "11000",
      "01010" when "11001",
      "01011" when "11010",
      "00000" when "11011",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(4 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
   instLUT: GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_28_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(4 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_9_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_28_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_20_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(4 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount281_out : std_logic_vector(4 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product34_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product34_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product316_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product316_8_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product316_8_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No27_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No108_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No28_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No109_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No29_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No30_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No111_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No31_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No112_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No32_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No5_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No113_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No33_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No105_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No6_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No34_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No35_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add11_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add11_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No241_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No18_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No36_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No19_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No37_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No20_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No38_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add3_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add3_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add3_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add3_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No111_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No112_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No113_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add12_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add12_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add12_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add12_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product11_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product11_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product11_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product11_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product21_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product21_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product21_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product21_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No90_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No91_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No93_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No94_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No95_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No42_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No33_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No233_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No125_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product12_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product12_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product22_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product22_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product6_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product6_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product23_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product23_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product33_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product33_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product33_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product33_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No18_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No19_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No20_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No21_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No22_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No23_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No24_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Subtract4_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Subtract4_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No25_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Subtract4_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Subtract4_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No26_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product34_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product34_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product34_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product34_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Product10_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Product10_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product28_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product28_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product42_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product42_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Product213_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Product213_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product213_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product213_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product313_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product313_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product316_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product316_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No19_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No2_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No20_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Subtract18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Subtract18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No3_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No21_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Subtract18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Subtract18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No4_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No22_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Subtract18_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Subtract18_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No5_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No23_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Subtract18_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Subtract18_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No6_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No24_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Subtract18_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Subtract18_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No7_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No25_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Subtract18_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Subtract18_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No8_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay45No26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Subtract22_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Subtract22_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Subtract22_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Subtract22_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Subtract22_7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Subtract22_7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Subtract22_8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Subtract22_8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount281_instance: ModuloCounter_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount281_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg115_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg125_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg135_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg145_out;
SharedReg155_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg165_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg175_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg145_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg185_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg198_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
SharedReg211_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg211_out;
SharedReg224_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg237_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg250_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg250_out;
SharedReg263_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg276_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg289_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg211_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg250_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg32_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg67_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg74_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg46_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg67_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg67_out;
SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg60_out;
SharedReg74_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg67_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg39_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg46_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg53_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg60_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg105_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg115_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg125_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg135_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg145_out;
SharedReg155_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg165_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg175_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg145_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg32_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg67_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg74_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg46_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg32_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg67_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg74_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg46_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg95_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg105_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg115_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg125_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg135_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg145_out;
SharedReg155_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg165_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg185_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg198_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
SharedReg211_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg211_out;
SharedReg224_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg237_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg250_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg250_out;
SharedReg263_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg276_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg289_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg211_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg250_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg67_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg74_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg46_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg115_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg125_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg135_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg145_out;
SharedReg155_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg165_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg175_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg145_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg185_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg198_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
SharedReg211_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg211_out;
SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg237_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg250_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg250_out;
SharedReg263_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg276_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg289_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg211_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg250_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg185_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg198_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
SharedReg211_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg211_out;
SharedReg224_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg237_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg250_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg250_out;
SharedReg263_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg276_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg289_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg211_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg250_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg32_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg39_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg46_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg53_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg60_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg67_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg74_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg81_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg88_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg46_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg105_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg115_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg125_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg135_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg145_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg145_out;
SharedReg155_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg165_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg175_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg175_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg125_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg145_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg185_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg198_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
SharedReg211_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg211_out;
SharedReg224_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg237_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg250_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg250_out;
SharedReg263_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg263_out;
SharedReg276_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg289_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg289_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg211_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg250_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg263_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg985_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg998_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg1011_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1011_out;
SharedReg1024_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1024_out;
SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1037_out;
SharedReg1050_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1050_out;
SharedReg1063_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg1076_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1076_out;
SharedReg1089_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1089_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1011_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1024_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1050_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1076_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1089_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg1142_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1150_out;
SharedReg1110_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1134_out;
SharedReg1158_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1142_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1150_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1110_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1118_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1126_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1134_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg1110_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg783_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg796_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg796_out;
SharedReg809_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg809_out;
SharedReg822_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg835_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg848_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg848_out;
SharedReg861_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg861_out;
SharedReg874_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg874_out;
SharedReg887_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg887_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg796_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg809_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg822_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg861_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg874_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg783_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg796_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg796_out;
SharedReg809_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg809_out;
SharedReg822_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg835_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg848_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg848_out;
SharedReg861_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg861_out;
SharedReg874_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg874_out;
SharedReg887_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg887_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg796_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg809_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg822_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg861_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg874_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg985_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg1011_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1011_out;
SharedReg1024_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1024_out;
SharedReg1037_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1037_out;
SharedReg1050_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1050_out;
SharedReg1063_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg1076_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1076_out;
SharedReg1089_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1089_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1011_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1024_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1037_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1050_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1076_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1089_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg1110_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg783_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg796_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg796_out;
SharedReg809_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg809_out;
SharedReg822_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg835_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg848_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg848_out;
SharedReg861_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg861_out;
SharedReg874_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg874_out;
SharedReg887_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg887_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg796_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg809_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg822_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg861_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg874_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg1110_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg511_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg511_out;
SharedReg525_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg525_out;
SharedReg539_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg539_out;
SharedReg553_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg553_out;
SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg567_out;
SharedReg581_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg581_out;
SharedReg595_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg595_out;
SharedReg609_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg609_out;
SharedReg623_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg623_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg511_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg525_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg539_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg553_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg581_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg595_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg609_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg623_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg985_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg998_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg1011_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1011_out;
SharedReg1024_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1024_out;
SharedReg1037_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1037_out;
SharedReg1050_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1050_out;
SharedReg1063_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg1076_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1076_out;
SharedReg1089_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1089_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1011_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1024_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1037_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1050_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1076_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1089_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg1110_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg985_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg1011_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1011_out;
SharedReg1024_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1024_out;
SharedReg1037_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1037_out;
SharedReg1050_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1050_out;
SharedReg1063_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg1076_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1076_out;
SharedReg1089_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1089_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1011_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1024_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1037_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1050_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1076_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1089_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg1110_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg985_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg1011_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1011_out;
SharedReg1024_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1024_out;
SharedReg1037_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1037_out;
SharedReg1050_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1050_out;
SharedReg1063_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg1076_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast <= SharedReg1076_out;
SharedReg1089_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast <= SharedReg1089_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1011_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1024_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1037_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1050_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1076_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1089_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg1110_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1118_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1126_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1134_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1142_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1142_out;
SharedReg1150_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1150_out;
SharedReg1158_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1166_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast <= SharedReg1166_out;
SharedReg1174_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1126_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1142_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1150_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1166_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg313_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg313_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg461_out;
SharedReg465_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg465_out;
SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg515_out;
SharedReg100_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg100_out;
SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg516_out;
SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg190_out;
SharedReg986_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg986_out;
SharedReg1112_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1112_out;
SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg305_out;
SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg515_out;
SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg515_out;
SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg99_out;
SharedReg194_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg194_out;
Delay8No27_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast <= Delay8No27_out;
SharedReg518_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg518_out;
SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg783_out;
SharedReg511_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg511_out;
SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg783_out;
SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg516_out;
SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg191_out;
SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg191_out;
SharedReg520_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg520_out;
SharedReg996_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg996_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg313_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg986_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1112_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg305_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg194_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay8No27_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg518_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg511_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg783_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg191_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg520_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg996_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg6_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg465_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg515_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg100_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg516_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

Delay27No_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= Delay27No_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg649_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg649_out;
Delay6No108_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= Delay6No108_out;
SharedReg519_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg519_out;
SharedReg193_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg193_out;
SharedReg521_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg104_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg104_out;
SharedReg1110_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
SharedReg985_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg985_out;
SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg303_out;
SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg785_out;
SharedReg513_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg513_out;
SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg303_out;
SharedReg197_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg197_out;
SharedReg410_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg410_out;
SharedReg788_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg788_out;
SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg511_out;
SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg785_out;
SharedReg1111_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1111_out;
SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg511_out;
SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg303_out;
SharedReg34_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg34_out;
SharedReg988_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg988_out;
SharedReg786_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg786_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay27No_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg104_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg985_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg513_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg197_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg410_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg788_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg785_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1111_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg511_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg303_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg34_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg988_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg786_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg649_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No108_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg519_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg193_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg204_out;
SharedReg534_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1009_out;
SharedReg325_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg325_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg467_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg467_out;
SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg471_out;
SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg529_out;
SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg110_out;
SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg530_out;
SharedReg203_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg203_out;
SharedReg999_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg999_out;
SharedReg1120_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1120_out;
SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg317_out;
SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg529_out;
SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg529_out;
SharedReg109_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg109_out;
SharedReg207_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg207_out;
Delay8No28_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast <= Delay8No28_out;
SharedReg532_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg532_out;
SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg796_out;
SharedReg525_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg525_out;
SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg796_out;
SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg530_out;
SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg204_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg110_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg203_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg999_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1120_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg317_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg529_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg109_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg207_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay8No28_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg532_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg525_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg796_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg530_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg204_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg325_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg6_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg467_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg41_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg1001_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg799_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg799_out;
Delay27No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= Delay27No1_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg654_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg654_out;
Delay6No109_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= Delay6No109_out;
SharedReg533_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg533_out;
SharedReg206_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg206_out;
SharedReg535_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg535_out;
SharedReg114_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg114_out;
SharedReg1118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1118_out;
SharedReg998_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg998_out;
SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg315_out;
SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg798_out;
SharedReg527_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg527_out;
SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg315_out;
SharedReg210_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg210_out;
SharedReg415_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg415_out;
SharedReg801_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg801_out;
SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg525_out;
SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg798_out;
SharedReg1119_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1119_out;
SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg525_out;
SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg315_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg533_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg206_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg535_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg114_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1118_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg998_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg527_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg799_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg210_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg415_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg801_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg798_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1119_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg525_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg315_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay27No1_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg654_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay6No109_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg809_out;
SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg544_out;
SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg217_out;
SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg217_out;
SharedReg548_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg1022_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1022_out;
SharedReg337_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg337_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg473_out;
SharedReg477_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg477_out;
SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg543_out;
SharedReg120_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg120_out;
SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg544_out;
SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg216_out;
SharedReg1012_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1012_out;
SharedReg1128_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1128_out;
SharedReg329_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg329_out;
SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg543_out;
SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg543_out;
SharedReg119_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg119_out;
SharedReg220_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg220_out;
Delay8No29_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast <= Delay8No29_out;
SharedReg546_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg546_out;
SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg809_out;
SharedReg539_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg539_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg477_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg120_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg544_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1012_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1128_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg329_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg543_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg119_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg220_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay8No29_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg546_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg809_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg539_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1022_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg337_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg6_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg1127_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1127_out;
SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg539_out;
SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg327_out;
SharedReg48_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg48_out;
SharedReg1014_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1014_out;
SharedReg812_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg812_out;
Delay27No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= Delay27No2_out;
SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg659_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg659_out;
Delay6No110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= Delay6No110_out;
SharedReg547_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg547_out;
SharedReg219_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg219_out;
SharedReg549_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg549_out;
SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg124_out;
SharedReg1126_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1126_out;
SharedReg1011_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1011_out;
SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg327_out;
SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg811_out;
SharedReg541_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg541_out;
SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg327_out;
SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg223_out;
SharedReg420_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg420_out;
SharedReg814_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg814_out;
SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg539_out;
SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg811_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1127_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg659_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay6No110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg547_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg219_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg549_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg124_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1126_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1011_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg541_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg223_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg420_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg814_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg539_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg811_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg48_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1014_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg812_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay27No2_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg822_out;
SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg558_out;
SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg230_out;
SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg230_out;
SharedReg562_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg1035_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1035_out;
SharedReg349_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg349_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
SharedReg479_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg479_out;
SharedReg483_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg483_out;
SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg557_out;
SharedReg130_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg130_out;
SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg558_out;
SharedReg229_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg229_out;
SharedReg1025_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1025_out;
SharedReg1136_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1136_out;
SharedReg341_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg341_out;
SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg557_out;
SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg557_out;
SharedReg129_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg129_out;
SharedReg233_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg233_out;
Delay8No30_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast <= Delay8No30_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg6_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg479_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg483_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg130_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg229_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg553_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1025_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1136_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg341_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg557_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg129_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg233_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay8No30_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg822_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg558_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg230_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1035_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg349_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg827_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg827_out;
SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg553_out;
SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg824_out;
SharedReg1135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1135_out;
SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg553_out;
SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg339_out;
SharedReg55_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg55_out;
SharedReg1027_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1027_out;
SharedReg825_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg825_out;
Delay27No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= Delay27No3_out;
SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
SharedReg664_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg664_out;
Delay6No111_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast <= Delay6No111_out;
SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg561_out;
SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg232_out;
SharedReg563_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg563_out;
SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg134_out;
SharedReg1134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1134_out;
SharedReg1024_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1024_out;
SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg339_out;
SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg824_out;
SharedReg555_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg555_out;
SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg339_out;
SharedReg236_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg236_out;
SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg425_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg827_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg664_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay6No111_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg563_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1024_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg824_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg555_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg236_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg425_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg553_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg339_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg55_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1027_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg825_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay27No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg139_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg139_out;
SharedReg246_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg246_out;
Delay8No31_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= Delay8No31_out;
SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg574_out;
SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg567_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg567_out;
SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg835_out;
SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg572_out;
SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg243_out;
SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg243_out;
SharedReg576_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg576_out;
SharedReg1048_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1048_out;
SharedReg361_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg361_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg12_out;
SharedReg485_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg485_out;
SharedReg489_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg489_out;
SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg571_out;
SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg140_out;
SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg572_out;
SharedReg242_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg242_out;
SharedReg1038_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1038_out;
SharedReg1144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1144_out;
SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg353_out;
SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg571_out;
SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg571_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg139_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg246_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg576_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1048_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg361_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg6_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg485_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg489_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay8No31_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg242_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1038_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg571_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg574_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg567_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg835_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg572_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg243_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg249_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg900_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg840_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg840_out;
SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg567_out;
SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg837_out;
SharedReg1143_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1143_out;
SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg351_out;
SharedReg62_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg1040_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1040_out;
SharedReg838_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg838_out;
Delay27No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= Delay27No4_out;
SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg28_out;
SharedReg669_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg669_out;
Delay6No112_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast <= Delay6No112_out;
SharedReg575_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg575_out;
SharedReg245_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg245_out;
SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg577_out;
SharedReg144_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg144_out;
SharedReg1142_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1142_out;
SharedReg1037_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1037_out;
SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg351_out;
SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg837_out;
SharedReg569_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg569_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1040_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg838_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay27No4_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg669_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay6No112_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg575_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg900_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg245_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg144_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1142_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1037_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg569_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg840_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg837_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1143_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg567_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg351_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_5_impl_out,
                 X => Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg365_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg365_out;
SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg585_out;
SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg585_out;
SharedReg149_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg149_out;
SharedReg259_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
Delay8No32_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast <= Delay8No32_out;
SharedReg588_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg588_out;
SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg848_out;
SharedReg581_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg581_out;
SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg848_out;
SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg586_out;
SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg256_out;
SharedReg590_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg590_out;
SharedReg1061_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1061_out;
SharedReg373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg373_out;
SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg12_out;
SharedReg491_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg491_out;
SharedReg495_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg495_out;
SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg585_out;
SharedReg150_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg150_out;
SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg586_out;
SharedReg255_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg255_out;
SharedReg1051_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1051_out;
SharedReg1152_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1152_out;
   MUX_Add2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg365_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg256_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg590_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1061_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg373_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg4_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg6_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg491_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg495_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg585_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg150_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg586_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg255_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1051_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1152_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg149_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay8No32_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg588_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg581_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_5_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_0_out,
                 Y => Delay1No42_out);

SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg363_out;
SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg850_out;
SharedReg583_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg583_out;
SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg363_out;
SharedReg262_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg453_out;
SharedReg853_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg853_out;
SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg581_out;
SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg1151_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1151_out;
SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg581_out;
SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg363_out;
SharedReg69_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg69_out;
SharedReg1053_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1053_out;
SharedReg851_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg851_out;
Delay27No5_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast <= Delay27No5_out;
SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg28_out;
SharedReg674_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg674_out;
Delay6No113_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast <= Delay6No113_out;
SharedReg589_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg589_out;
SharedReg258_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg258_out;
SharedReg591_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg591_out;
SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg154_out;
SharedReg1150_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1150_out;
SharedReg1050_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1050_out;
   MUX_Add2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg69_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1053_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg851_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay27No5_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg22_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg583_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg674_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay6No113_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg589_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg258_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg591_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg154_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1150_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1050_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg363_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg453_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg853_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg581_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1151_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_5_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_6_impl_out,
                 X => Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg268_out;
SharedReg1064_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1064_out;
SharedReg1160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1160_out;
SharedReg377_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg377_out;
SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg599_out;
SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg599_out;
SharedReg159_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg159_out;
SharedReg272_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg272_out;
Delay8No33_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast <= Delay8No33_out;
SharedReg602_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg602_out;
SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg861_out;
SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg595_out;
SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg861_out;
SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg600_out;
SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg269_out;
SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg269_out;
SharedReg604_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg604_out;
SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1074_out;
SharedReg385_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg385_out;
SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg12_out;
SharedReg679_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg679_out;
Delay6No105_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast <= Delay6No105_out;
SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg599_out;
SharedReg160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg160_out;
SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg600_out;
   MUX_Add2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg268_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1064_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg861_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg269_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg604_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1074_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg385_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg4_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg679_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay6No105_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg160_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg377_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg599_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg159_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg272_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay8No33_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg602_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_6_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_0_out,
                 Y => Delay1No44_out);

SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg1158_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1158_out;
SharedReg1063_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1063_out;
SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg375_out;
SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg863_out;
SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg597_out;
SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg375_out;
SharedReg275_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg275_out;
SharedReg440_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg440_out;
SharedReg866_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg866_out;
SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg595_out;
SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg863_out;
SharedReg1159_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1159_out;
SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg595_out;
SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg375_out;
SharedReg76_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg76_out;
SharedReg1066_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1066_out;
SharedReg864_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg864_out;
Delay27No6_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast <= Delay27No6_out;
SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg28_out;
SharedReg767_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg767_out;
SharedReg771_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg771_out;
SharedReg603_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg603_out;
SharedReg271_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg271_out;
SharedReg605_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg605_out;
   MUX_Add2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1158_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1159_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg76_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1066_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg864_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay27No6_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1063_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg20_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg22_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg767_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg771_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg603_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg271_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg605_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg863_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg375_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg275_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg440_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg866_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_6_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add2_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_7_impl_out,
                 X => Delay1No46_out_to_Add2_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add2_7_impl_parent_implementedSystem_port_1_cast);

SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg613_out;
SharedReg170_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg614_out;
SharedReg281_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg281_out;
SharedReg1077_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1077_out;
SharedReg1168_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1168_out;
SharedReg389_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg389_out;
SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg613_out;
SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg613_out;
SharedReg169_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg169_out;
SharedReg285_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg285_out;
Delay8No34_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast <= Delay8No34_out;
SharedReg616_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg616_out;
SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg874_out;
SharedReg609_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg609_out;
SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg874_out;
SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg614_out;
SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg282_out;
SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg282_out;
SharedReg618_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg618_out;
SharedReg1087_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1087_out;
SharedReg397_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg397_out;
SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg12_out;
SharedReg684_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg684_out;
SharedReg688_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg688_out;
   MUX_Add2_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg285_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay8No34_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg616_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg609_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg874_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg282_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg618_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg614_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1087_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg397_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg4_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg6_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg12_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg684_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg688_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg281_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1077_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1168_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg389_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg613_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg169_out_to_MUX_Add2_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_7_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_7_impl_0_out,
                 Y => Delay1No46_out);

SharedReg617_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg617_out;
SharedReg284_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg284_out;
SharedReg619_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg619_out;
SharedReg174_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg174_out;
SharedReg1166_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1166_out;
SharedReg1076_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1076_out;
SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg387_out;
SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg876_out;
SharedReg611_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg611_out;
SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg387_out;
SharedReg288_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg288_out;
SharedReg502_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg502_out;
SharedReg879_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg879_out;
SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg609_out;
SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg876_out;
SharedReg1167_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1167_out;
SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg609_out;
SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg387_out;
SharedReg83_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg83_out;
SharedReg1079_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1079_out;
SharedReg877_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg877_out;
Delay27No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast <= Delay27No7_out;
SharedReg16_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg28_out;
SharedReg773_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg773_out;
SharedReg777_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg777_out;
   MUX_Add2_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg617_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg284_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg288_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg502_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg879_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1167_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg609_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg83_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1079_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg619_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg877_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay27No7_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg16_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg20_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg22_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg28_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg773_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg777_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg174_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1166_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1076_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg876_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg611_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg387_out_to_MUX_Add2_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_7_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_7_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add2_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_8_impl_out,
                 X => Delay1No48_out_to_Add2_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add2_8_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg506_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg506_out;
SharedReg694_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg694_out;
SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg180_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg180_out;
SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg628_out;
SharedReg294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg294_out;
SharedReg1090_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1090_out;
SharedReg1176_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1176_out;
SharedReg401_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg401_out;
SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg627_out;
SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg627_out;
SharedReg179_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg179_out;
SharedReg298_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg298_out;
Delay8No35_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast <= Delay8No35_out;
SharedReg630_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg630_out;
SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg887_out;
SharedReg623_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg623_out;
SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg887_out;
SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg628_out;
SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg295_out;
SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg295_out;
SharedReg632_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg632_out;
SharedReg1100_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1100_out;
SharedReg409_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg409_out;
SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg4_out;
   MUX_Add2_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg401_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg179_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg298_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay8No35_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg630_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg623_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg887_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg506_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg295_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg632_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1100_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg409_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg4_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg694_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg180_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg628_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg294_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1090_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1176_out_to_MUX_Add2_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_8_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_8_impl_0_out,
                 Y => Delay1No48_out);

SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg28_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg690_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg690_out;
SharedReg731_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg731_out;
SharedReg631_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg631_out;
SharedReg297_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
SharedReg633_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg633_out;
SharedReg184_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg184_out;
SharedReg1174_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
SharedReg1089_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1089_out;
SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg399_out;
SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg889_out;
SharedReg625_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg625_out;
SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg399_out;
SharedReg301_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg301_out;
SharedReg637_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg637_out;
SharedReg892_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg892_out;
SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg623_out;
SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg889_out;
SharedReg1175_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1175_out;
SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg623_out;
SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg399_out;
SharedReg90_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg90_out;
SharedReg1092_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1092_out;
SharedReg890_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg890_out;
Delay27No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast <= Delay27No8_out;
SharedReg16_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg20_out;
   MUX_Add2_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg625_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg301_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg637_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg892_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg889_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1175_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg690_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg623_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg399_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg90_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1092_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg890_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay27No8_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg16_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg20_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg731_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg631_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg297_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg633_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg184_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1089_out_to_MUX_Add2_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add2_8_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_8_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No50_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg412_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg412_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg462_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg462_out;
SharedReg464_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg410_out;
SharedReg788_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg788_out;
SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg307_out;
SharedReg789_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg789_out;
SharedReg784_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg784_out;
SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg410_out;
SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg36_out;
SharedReg512_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg512_out;
SharedReg792_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg792_out;
SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg410_out;
SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg735_out;
SharedReg522_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg522_out;
SharedReg304_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg304_out;
SharedReg302_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg302_out;
SharedReg185_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg185_out;
SharedReg100_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg100_out;
SharedReg649_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg649_out;
SharedReg790_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg790_out;
SharedReg650_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg650_out;
SharedReg195_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg195_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg412_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg789_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg784_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg512_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg792_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg522_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg5_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg304_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg302_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg185_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg100_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg649_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg790_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg650_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg195_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg9_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg462_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg410_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg788_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg307_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No50_out);

SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg460_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg650_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg650_out;
SharedReg652_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg652_out;
SharedReg461_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg461_out;
SharedReg992_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg992_out;
SharedReg309_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg309_out;
SharedReg793_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg793_out;
SharedReg783_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg783_out;
SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg460_out;
SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg463_out;
SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg187_out;
SharedReg986_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg986_out;
SharedReg524_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg524_out;
SharedReg651_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg651_out;
SharedReg648_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg648_out;
SharedReg523_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg523_out;
SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg302_out;
SharedReg304_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg304_out;
SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg302_out;
SharedReg95_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg95_out;
SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg462_out;
SharedReg512_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg512_out;
SharedReg696_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg696_out;
SharedReg305_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg305_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg793_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg783_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg460_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg187_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg986_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg524_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg651_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg648_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg523_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg304_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg302_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg95_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg512_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg696_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg305_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg25_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg650_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg652_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg461_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg992_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg309_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No52_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg803_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg655_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg655_out;
SharedReg208_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg208_out;
SharedReg1104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1104_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg468_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg468_out;
SharedReg470_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg470_out;
SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg415_out;
SharedReg801_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg319_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg319_out;
SharedReg802_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg802_out;
SharedReg797_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg797_out;
SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg415_out;
SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg415_out;
SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg43_out;
SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg526_out;
SharedReg805_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg805_out;
SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg415_out;
SharedReg740_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg740_out;
SharedReg536_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg536_out;
SharedReg316_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg316_out;
SharedReg314_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg314_out;
SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg198_out;
SharedReg110_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg110_out;
SharedReg654_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg654_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg655_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg319_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg802_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg797_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg43_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg526_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg805_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg208_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg415_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg740_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg536_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg316_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg314_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg110_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg654_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg9_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg468_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg470_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No52_out);

SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg526_out;
SharedReg654_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg654_out;
SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg415_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg415_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg655_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg655_out;
SharedReg657_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg657_out;
SharedReg467_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg467_out;
SharedReg1005_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1005_out;
SharedReg321_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg321_out;
SharedReg806_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg806_out;
SharedReg796_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg796_out;
SharedReg466_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg466_out;
SharedReg469_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg469_out;
SharedReg200_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg200_out;
SharedReg999_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg999_out;
SharedReg538_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg538_out;
SharedReg656_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg656_out;
SharedReg653_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg653_out;
SharedReg537_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg537_out;
SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg314_out;
SharedReg316_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg316_out;
SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg314_out;
SharedReg105_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg105_out;
SharedReg468_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg468_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg526_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg654_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg467_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1005_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg321_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg806_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg796_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg466_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg469_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg200_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg999_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg538_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg317_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg656_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg653_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg537_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg316_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg314_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg105_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg468_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg415_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg25_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg655_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg657_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No54_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg211_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg120_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg120_out;
SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg473_out;
SharedReg816_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg474_out;
SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg221_out;
SharedReg1108_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1108_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg474_out;
SharedReg476_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg476_out;
SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg420_out;
SharedReg814_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg814_out;
SharedReg331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg331_out;
SharedReg815_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg815_out;
SharedReg810_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg810_out;
SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg420_out;
SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg420_out;
SharedReg50_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg50_out;
SharedReg540_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg540_out;
SharedReg818_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg818_out;
SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg420_out;
SharedReg745_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg745_out;
SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg550_out;
SharedReg328_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg328_out;
SharedReg326_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg326_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg476_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg814_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg331_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg815_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg810_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg50_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg540_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg818_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg745_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg328_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg326_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg816_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg474_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1108_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No54_out);

SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg115_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg115_out;
SharedReg422_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg422_out;
SharedReg540_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg540_out;
SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg473_out;
SharedReg329_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg329_out;
SharedReg420_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg420_out;
SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg660_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg660_out;
SharedReg662_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg662_out;
SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg473_out;
SharedReg1018_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1018_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg333_out;
SharedReg819_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg819_out;
SharedReg809_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg809_out;
SharedReg472_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg472_out;
SharedReg475_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg475_out;
SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg213_out;
SharedReg1012_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1012_out;
SharedReg552_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg552_out;
SharedReg661_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg661_out;
SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg658_out;
SharedReg551_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg551_out;
SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg326_out;
SharedReg328_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg328_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg115_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg660_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg662_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1018_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg819_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg809_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg472_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg475_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg422_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1012_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg552_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg661_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg551_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg328_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg540_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg473_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg329_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg420_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No56_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg564_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg564_out;
SharedReg340_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg340_out;
SharedReg338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg224_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg130_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
SharedReg479_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg479_out;
SharedReg829_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg480_out;
SharedReg234_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg234_out;
SharedReg911_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg911_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg7_out;
SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg480_out;
SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg482_out;
SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg425_out;
SharedReg827_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg827_out;
SharedReg343_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg343_out;
SharedReg828_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg828_out;
SharedReg823_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg823_out;
SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg425_out;
SharedReg57_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg57_out;
SharedReg554_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg554_out;
SharedReg831_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg831_out;
SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg425_out;
SharedReg750_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg750_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg564_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg9_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg482_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg827_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg343_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg828_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg338_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg823_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg57_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg554_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg831_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg425_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg750_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg224_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg479_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg480_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg234_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg911_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No56_out);

SharedReg565_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg340_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg340_out;
SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg338_out;
SharedReg125_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg125_out;
SharedReg911_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg911_out;
SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg479_out;
SharedReg341_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg341_out;
SharedReg425_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg425_out;
SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg23_out;
SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg665_out;
SharedReg667_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg667_out;
SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg479_out;
SharedReg1031_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1031_out;
SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg345_out;
SharedReg832_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg832_out;
SharedReg822_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg822_out;
SharedReg478_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg478_out;
SharedReg481_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg481_out;
SharedReg226_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg226_out;
SharedReg1025_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1025_out;
SharedReg566_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg566_out;
SharedReg666_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg666_out;
SharedReg663_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg663_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg667_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1031_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg832_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg340_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg822_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg478_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg481_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg226_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1025_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg566_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg666_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg663_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg338_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg125_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg911_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg479_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg341_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg425_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No58_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg844_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg844_out;
SharedReg900_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg756_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg578_out;
SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg350_out;
SharedReg237_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg237_out;
SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg140_out;
SharedReg485_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg485_out;
SharedReg842_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg842_out;
SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg486_out;
SharedReg247_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg247_out;
SharedReg902_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg902_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg7_out;
SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg486_out;
SharedReg488_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg488_out;
SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg430_out;
SharedReg840_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg840_out;
SharedReg355_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg355_out;
SharedReg841_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg841_out;
SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg836_out;
SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg430_out;
SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg430_out;
SharedReg64_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg64_out;
SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg568_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg844_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg247_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg902_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg9_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg7_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg486_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg488_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg756_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg840_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg355_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg841_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg430_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg64_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg568_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg237_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg485_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg842_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No58_out);

SharedReg580_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg580_out;
SharedReg671_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg671_out;
SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg484_out;
SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg579_out;
SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg350_out;
SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg352_out;
SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg350_out;
SharedReg135_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg135_out;
SharedReg902_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg902_out;
SharedReg568_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg485_out;
SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg353_out;
SharedReg430_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg430_out;
SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg23_out;
SharedReg670_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg670_out;
SharedReg672_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg672_out;
SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg485_out;
SharedReg1044_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1044_out;
SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg357_out;
SharedReg845_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg845_out;
SharedReg835_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg835_out;
SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg484_out;
SharedReg487_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg487_out;
SharedReg239_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg239_out;
SharedReg1038_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1038_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg580_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg671_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg353_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg430_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg25_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg670_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg672_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg485_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1044_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg357_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg845_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg835_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg484_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg487_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg239_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1038_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg350_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg135_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg902_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add11_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_5_impl_out,
                 X => Delay1No60_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast);

SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg453_out;
SharedReg71_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg582_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg582_out;
SharedReg857_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg857_out;
SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg453_out;
SharedReg762_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg762_out;
SharedReg592_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg592_out;
SharedReg364_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg364_out;
SharedReg362_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg362_out;
SharedReg250_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg250_out;
SharedReg150_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg150_out;
SharedReg491_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg491_out;
SharedReg855_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg855_out;
SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg492_out;
SharedReg260_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg260_out;
SharedReg455_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg455_out;
SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg7_out;
SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg492_out;
SharedReg494_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg494_out;
SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg435_out;
SharedReg853_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg853_out;
SharedReg367_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg367_out;
SharedReg854_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg854_out;
SharedReg849_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg849_out;
SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg435_out;
   MUX_Add11_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg150_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg491_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg855_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg260_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg455_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg9_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg582_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg492_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg494_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg853_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg367_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg854_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg849_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg435_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg857_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg453_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg762_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg592_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg364_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg362_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg250_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_5_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_0_out,
                 Y => Delay1No60_out);

SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg493_out;
SharedReg252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg1051_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1051_out;
SharedReg594_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg594_out;
SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg493_out;
SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg490_out;
SharedReg593_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg593_out;
SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg364_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg364_out;
SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg362_out;
SharedReg145_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg145_out;
SharedReg455_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg455_out;
SharedReg582_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg582_out;
SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg491_out;
SharedReg365_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg365_out;
SharedReg435_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg435_out;
SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg23_out;
SharedReg675_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg675_out;
SharedReg677_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg677_out;
SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg491_out;
SharedReg1057_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1057_out;
SharedReg369_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg369_out;
SharedReg858_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg858_out;
SharedReg848_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg848_out;
SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg490_out;
   MUX_Add11_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg145_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg455_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg582_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg365_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg435_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg21_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg25_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1051_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg675_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg677_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg491_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1057_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg369_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg858_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg848_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg594_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg493_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg490_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg593_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg364_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg362_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_5_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add11_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_6_impl_out,
                 X => Delay1No62_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast);

SharedReg867_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg867_out;
SharedReg862_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg440_out;
SharedReg456_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg456_out;
SharedReg78_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg78_out;
SharedReg596_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg596_out;
SharedReg870_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg870_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg440_out;
SharedReg923_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg923_out;
SharedReg606_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg606_out;
SharedReg376_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg374_out;
SharedReg263_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg263_out;
SharedReg160_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg160_out;
SharedReg679_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg679_out;
SharedReg868_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg868_out;
SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg680_out;
SharedReg273_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg273_out;
SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg442_out;
SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg7_out;
SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg680_out;
SharedReg682_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg682_out;
SharedReg496_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg496_out;
SharedReg866_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg866_out;
SharedReg379_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg379_out;
   MUX_Add11_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg867_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg376_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg374_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg263_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg160_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg679_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg868_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg273_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg5_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg9_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg7_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg680_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg682_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg496_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg866_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg379_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg456_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg78_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg596_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg870_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg923_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg606_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_6_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_0_out,
                 Y => Delay1No62_out);

SharedReg871_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg861_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg861_out;
SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg496_out;
SharedReg499_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg499_out;
SharedReg265_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg1064_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1064_out;
SharedReg608_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg608_out;
SharedReg681_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg681_out;
SharedReg678_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg678_out;
SharedReg607_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg607_out;
SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg376_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg374_out;
SharedReg155_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg155_out;
SharedReg442_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg442_out;
SharedReg596_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg596_out;
SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg679_out;
SharedReg377_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg377_out;
SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg496_out;
SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg23_out;
SharedReg768_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg768_out;
SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg770_out;
SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg679_out;
SharedReg1070_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1070_out;
SharedReg381_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg381_out;
   MUX_Add11_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg861_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg376_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg374_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg155_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg442_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg596_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg377_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg496_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg21_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg25_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg23_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg768_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg679_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1070_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg381_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg499_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1064_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg608_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg681_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg678_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg607_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_6_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add11_7_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add11_7_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add11_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_7_impl_out,
                 X => Delay1No64_out_to_Add11_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add11_7_impl_parent_implementedSystem_port_1_cast);

SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg502_out;
SharedReg879_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg879_out;
SharedReg391_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg880_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg880_out;
SharedReg875_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg875_out;
SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg502_out;
SharedReg444_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg444_out;
SharedReg85_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg85_out;
SharedReg610_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg610_out;
SharedReg883_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg883_out;
SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg502_out;
SharedReg929_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg929_out;
SharedReg620_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg620_out;
SharedReg388_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg388_out;
SharedReg386_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg386_out;
SharedReg276_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg276_out;
SharedReg170_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg170_out;
SharedReg684_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg684_out;
SharedReg881_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg881_out;
SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg685_out;
SharedReg286_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg286_out;
SharedReg504_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg504_out;
SharedReg1_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg7_out;
SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg685_out;
SharedReg687_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg687_out;
   MUX_Add11_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg879_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg929_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg620_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg388_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg386_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg276_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg170_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg684_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg881_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg391_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg286_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg504_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg5_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg9_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg7_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg685_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg687_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg880_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg875_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg502_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg444_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg85_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg610_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg883_out_to_MUX_Add11_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_7_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_7_impl_0_out,
                 Y => Delay1No64_out);

SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg684_out;
SharedReg1083_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1083_out;
SharedReg393_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg393_out;
SharedReg884_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg884_out;
SharedReg874_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg874_out;
SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg642_out;
Delay4No241_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_7_cast <= Delay4No241_out;
SharedReg278_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg278_out;
SharedReg1077_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1077_out;
SharedReg622_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg622_out;
SharedReg686_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg686_out;
SharedReg683_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg683_out;
SharedReg621_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg621_out;
SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg386_out;
SharedReg388_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg388_out;
SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg386_out;
SharedReg165_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg165_out;
SharedReg504_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg504_out;
SharedReg610_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg610_out;
SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg684_out;
SharedReg389_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg389_out;
SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg642_out;
SharedReg17_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg23_out;
SharedReg774_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg774_out;
SharedReg776_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg776_out;
   MUX_Add11_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1083_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg686_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg683_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg621_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg388_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg386_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg165_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg504_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg610_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg684_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg393_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg389_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg17_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg21_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg25_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg23_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg774_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg776_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg884_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg874_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg642_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay4No241_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg278_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1077_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg622_out_to_MUX_Add11_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_7_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_7_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add11_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_8_impl_out,
                 X => Delay1No66_out_to_Add11_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add11_8_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg7_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg507_out;
SharedReg693_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg693_out;
SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg450_out;
SharedReg892_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg892_out;
SharedReg403_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg403_out;
SharedReg893_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg893_out;
SharedReg888_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg888_out;
SharedReg637_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg637_out;
SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg450_out;
SharedReg92_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg92_out;
SharedReg624_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg624_out;
SharedReg896_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg896_out;
SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg450_out;
SharedReg729_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg729_out;
SharedReg634_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg634_out;
SharedReg400_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg400_out;
SharedReg398_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg398_out;
SharedReg289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg289_out;
SharedReg180_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg180_out;
SharedReg690_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg690_out;
SharedReg894_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg894_out;
SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg507_out;
SharedReg299_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg299_out;
SharedReg452_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg452_out;
SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg5_out;
   MUX_Add11_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg92_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg624_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg896_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg729_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg634_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg400_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg398_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg289_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg180_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg690_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg894_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg507_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg299_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg452_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg5_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg693_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg450_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg892_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg403_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg893_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg888_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg637_out_to_MUX_Add11_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_8_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_8_impl_0_out,
                 Y => Delay1No66_out);

SharedReg25_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg23_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg691_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg691_out;
SharedReg730_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg730_out;
SharedReg451_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg451_out;
SharedReg1096_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1096_out;
SharedReg405_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg405_out;
SharedReg897_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg897_out;
SharedReg887_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg887_out;
SharedReg450_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg450_out;
SharedReg508_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg508_out;
SharedReg291_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg291_out;
SharedReg1090_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1090_out;
SharedReg636_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg636_out;
SharedReg692_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg692_out;
SharedReg505_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg505_out;
SharedReg635_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg635_out;
SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg398_out;
SharedReg400_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg400_out;
SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg398_out;
SharedReg175_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg175_out;
SharedReg507_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg507_out;
SharedReg624_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg624_out;
SharedReg727_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg727_out;
SharedReg401_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg401_out;
SharedReg689_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg689_out;
SharedReg17_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg21_out;
   MUX_Add11_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg508_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg291_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1090_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg636_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg692_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg505_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg635_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg400_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg398_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg691_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg175_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg507_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg624_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg727_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg401_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg689_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg17_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg21_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg730_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg451_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1096_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg405_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg897_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg450_out_to_MUX_Add11_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add11_8_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_8_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_0_impl_out,
                 X => Delay1No68_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg410_out;
SharedReg695_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg695_out;
SharedReg650_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg650_out;
SharedReg189_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg189_out;
Delay9No18_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast <= Delay9No18_out;
SharedReg307_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg307_out;
SharedReg96_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg96_out;
SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg733_out;
SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg412_out;
SharedReg35_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg35_out;
SharedReg186_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg186_out;
SharedReg993_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg993_out;
SharedReg648_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg648_out;
SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg733_out;
SharedReg102_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg102_out;
SharedReg1116_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1116_out;
SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg410_out;
SharedReg518_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg518_out;
SharedReg515_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg515_out;
SharedReg696_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg696_out;
SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg412_out;
SharedReg940_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg940_out;
SharedReg460_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg460_out;
   MUX_Add3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg307_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg96_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg35_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg186_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg993_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg648_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg733_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg102_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg13_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1116_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg518_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg515_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg696_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg412_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg940_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg460_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg10_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg410_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg695_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg650_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg189_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay9No18_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_0_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_0_out,
                 Y => Delay1No68_out);

SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg940_out;
SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg941_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg941_out;
SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg732_out;
SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg695_out;
SharedReg308_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg648_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg648_out;
SharedReg309_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg309_out;
SharedReg95_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg939_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg939_out;
SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg695_out;
SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg303_out;
SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg303_out;
SharedReg795_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg795_out;
SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg940_out;
SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg732_out;
SharedReg196_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg196_out;
SharedReg794_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg794_out;
SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg461_out;
SharedReg511_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg511_out;
SharedReg783_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg783_out;
SharedReg734_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg734_out;
SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg461_out;
SharedReg1103_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1103_out;
Delay9No36_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_28_cast <= Delay9No36_out;
   MUX_Add3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg309_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg939_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg303_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg795_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg940_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg196_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg29_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg794_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg511_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg783_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg734_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg461_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1103_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay9No36_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg26_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg941_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg732_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg695_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg648_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_0_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_1_impl_out,
                 X => Delay1No70_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg417_out;
SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg738_out;
SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg702_out;
SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg415_out;
SharedReg701_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg701_out;
SharedReg655_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg655_out;
SharedReg202_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg202_out;
Delay9No19_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast <= Delay9No19_out;
SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg319_out;
SharedReg106_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg106_out;
SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg738_out;
SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg417_out;
SharedReg42_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg42_out;
SharedReg199_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg199_out;
SharedReg1006_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1006_out;
SharedReg653_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg653_out;
SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg738_out;
SharedReg112_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg112_out;
SharedReg1124_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1124_out;
SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg415_out;
SharedReg532_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg532_out;
SharedReg529_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg529_out;
SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg702_out;
   MUX_Add3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg655_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay9No19_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg106_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg417_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg42_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg199_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1006_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg653_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg738_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg112_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1124_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg532_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg529_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg702_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg10_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg415_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg701_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_1_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_0_out,
                 Y => Delay1No70_out);

SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg467_out;
SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg947_out;
Delay9No37_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast <= Delay9No37_out;
SharedReg738_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg738_out;
SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg948_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg948_out;
SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg737_out;
SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg701_out;
SharedReg320_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg320_out;
SharedReg653_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg653_out;
SharedReg321_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg321_out;
SharedReg105_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg105_out;
SharedReg946_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg946_out;
SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg701_out;
SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg315_out;
SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg315_out;
SharedReg808_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg808_out;
SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg947_out;
SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg737_out;
SharedReg209_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg209_out;
SharedReg807_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg807_out;
SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg467_out;
SharedReg525_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg525_out;
SharedReg796_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg796_out;
SharedReg739_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg739_out;
   MUX_Add3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg320_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg653_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg321_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg105_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg946_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg701_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg315_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg808_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay9No37_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg947_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg209_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg807_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg467_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg525_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg796_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg739_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg738_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg26_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg948_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg737_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_1_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_2_impl_out,
                 X => Delay1No72_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg546_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg546_out;
SharedReg543_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg543_out;
SharedReg659_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg659_out;
SharedReg1108_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1108_out;
SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg708_out;
SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg420_out;
SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg708_out;
SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg420_out;
SharedReg707_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg707_out;
SharedReg660_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg660_out;
SharedReg215_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg215_out;
Delay9No20_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_16_cast <= Delay9No20_out;
SharedReg331_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg331_out;
SharedReg116_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg116_out;
SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg743_out;
SharedReg422_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg422_out;
SharedReg49_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg49_out;
SharedReg212_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg212_out;
SharedReg1019_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1019_out;
SharedReg658_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg658_out;
SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg743_out;
SharedReg122_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg122_out;
SharedReg1132_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1132_out;
SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg420_out;
   MUX_Add3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg546_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg543_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg707_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg660_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg215_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay9No20_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg331_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg116_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg422_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg659_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg49_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg212_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1019_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg658_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg743_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg122_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1132_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1108_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg420_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg708_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg10_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_2_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_0_out,
                 Y => Delay1No72_out);

SharedReg539_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg539_out;
SharedReg809_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg809_out;
SharedReg709_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg709_out;
SharedReg421_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg421_out;
SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg743_out;
Delay9No38_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast <= Delay9No38_out;
SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg743_out;
SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg955_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg955_out;
SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg742_out;
SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg707_out;
SharedReg332_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg332_out;
SharedReg658_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg658_out;
SharedReg333_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg333_out;
SharedReg115_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg115_out;
SharedReg953_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg953_out;
SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg707_out;
SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg327_out;
SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg327_out;
SharedReg821_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg821_out;
SharedReg954_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg954_out;
SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg742_out;
SharedReg222_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg222_out;
SharedReg820_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg820_out;
SharedReg473_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg473_out;
   MUX_Add3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg539_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg809_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg955_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg332_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg658_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg333_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg115_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg953_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg707_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg709_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg327_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg821_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg954_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg742_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg222_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg820_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg473_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg421_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay9No38_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg743_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg26_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_2_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_3_impl_out,
                 X => Delay1No74_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg132_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg1140_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1140_out;
SharedReg909_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg560_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg560_out;
SharedReg557_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg557_out;
SharedReg664_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg664_out;
SharedReg911_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg911_out;
SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg714_out;
SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg425_out;
SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg714_out;
SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg8_out;
SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg425_out;
SharedReg713_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg713_out;
SharedReg665_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg665_out;
SharedReg228_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg228_out;
SharedReg752_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg752_out;
SharedReg343_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg343_out;
SharedReg126_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg126_out;
SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg748_out;
SharedReg427_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg427_out;
SharedReg56_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg56_out;
SharedReg225_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg225_out;
SharedReg1032_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1032_out;
SharedReg663_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg663_out;
SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg748_out;
   MUX_Add3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1140_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg13_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg10_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg8_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg713_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg665_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg228_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg752_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg343_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg909_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg126_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg427_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg56_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg225_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1032_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg663_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg748_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg560_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg557_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg664_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg911_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg425_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg714_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_3_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_0_out,
                 Y => Delay1No74_out);

SharedReg235_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg833_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg833_out;
SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg553_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg553_out;
SharedReg822_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg822_out;
SharedReg665_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg665_out;
SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg748_out;
SharedReg919_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg919_out;
SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg748_out;
SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
SharedReg915_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg915_out;
SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg747_out;
SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg713_out;
SharedReg344_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg344_out;
SharedReg663_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg663_out;
SharedReg345_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg345_out;
SharedReg125_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg125_out;
SharedReg913_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg913_out;
SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg713_out;
SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg339_out;
SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg339_out;
SharedReg834_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg834_out;
SharedReg914_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg914_out;
SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg747_out;
   MUX_Add3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg833_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg29_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg26_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg915_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg344_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg663_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg345_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg125_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg913_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg713_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg339_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg834_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg914_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg747_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg553_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg822_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg665_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg426_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg919_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg748_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_3_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_4_impl_out,
                 X => Delay1No76_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1045_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1045_out;
SharedReg484_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg484_out;
SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg720_out;
SharedReg142_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg142_out;
SharedReg1148_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1148_out;
SharedReg900_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg900_out;
SharedReg574_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg574_out;
SharedReg571_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg571_out;
SharedReg669_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg669_out;
SharedReg902_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg902_out;
SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg720_out;
SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg430_out;
SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg720_out;
SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg8_out;
SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg430_out;
SharedReg719_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg719_out;
SharedReg670_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg670_out;
SharedReg241_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg241_out;
SharedReg758_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg758_out;
SharedReg355_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg355_out;
SharedReg136_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg136_out;
SharedReg754_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg754_out;
SharedReg432_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg432_out;
SharedReg63_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg63_out;
SharedReg238_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg238_out;
   MUX_Add3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1045_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg484_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg13_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg10_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg8_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg430_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg719_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg670_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg720_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg241_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg758_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg355_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg136_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg754_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg432_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg63_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg238_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg142_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1148_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg900_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg574_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg571_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg669_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg902_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_4_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_0_out,
                 Y => Delay1No76_out);

SharedReg847_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg847_out;
SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg754_out;
SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg248_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg248_out;
SharedReg846_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg846_out;
SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg431_out;
SharedReg567_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg835_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg670_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg670_out;
SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg431_out;
SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg754_out;
SharedReg758_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg758_out;
SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg754_out;
SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg24_out;
SharedReg905_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg905_out;
SharedReg753_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg753_out;
SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg719_out;
SharedReg356_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg356_out;
SharedReg668_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg668_out;
SharedReg357_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg357_out;
SharedReg135_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg135_out;
SharedReg903_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg903_out;
SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg719_out;
SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg351_out;
SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg351_out;
   MUX_Add3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg847_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg754_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg29_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg24_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg905_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg753_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg356_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg668_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg357_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg135_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg903_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg719_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg351_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg248_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg846_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg670_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg431_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_4_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add3_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_5_impl_out,
                 X => Delay1No78_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast);

SharedReg437_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg437_out;
SharedReg70_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg70_out;
SharedReg251_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg251_out;
SharedReg1058_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1058_out;
SharedReg490_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg490_out;
SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg760_out;
SharedReg152_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg152_out;
SharedReg1156_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1156_out;
SharedReg453_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg453_out;
SharedReg588_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg588_out;
SharedReg585_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg585_out;
SharedReg674_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg674_out;
SharedReg455_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg455_out;
SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg760_out;
SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg435_out;
SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg760_out;
SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg8_out;
SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg435_out;
SharedReg759_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg759_out;
SharedReg675_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg675_out;
SharedReg254_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg254_out;
SharedReg938_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg938_out;
SharedReg367_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg367_out;
SharedReg146_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg146_out;
SharedReg933_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg933_out;
   MUX_Add3_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg437_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg70_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg585_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg674_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg455_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg13_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg10_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg251_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg435_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg759_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg675_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg254_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg938_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg367_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg146_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg933_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1058_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg490_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg760_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg152_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1156_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg453_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg588_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_5_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_5_impl_0_out,
                 Y => Delay1No78_out);

SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg363_out;
SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg363_out;
SharedReg860_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg860_out;
SharedReg760_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg760_out;
SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg759_out;
SharedReg261_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg859_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg859_out;
SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg436_out;
SharedReg581_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg581_out;
SharedReg848_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg848_out;
SharedReg675_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg675_out;
SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg436_out;
SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg933_out;
SharedReg938_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg938_out;
SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg933_out;
SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg24_out;
SharedReg458_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg458_out;
SharedReg932_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg932_out;
SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg759_out;
SharedReg368_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg368_out;
SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg673_out;
SharedReg369_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg369_out;
SharedReg145_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg145_out;
SharedReg456_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg456_out;
   MUX_Add3_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg848_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg675_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg938_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg933_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg29_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg26_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg363_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg458_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg932_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg368_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg673_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg369_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg145_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg456_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg860_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg760_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg759_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg859_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg436_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg581_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_5_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_5_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add3_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_6_impl_out,
                 X => Delay1No80_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast);

SharedReg379_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg156_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg921_out;
SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg442_out;
SharedReg77_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg264_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg264_out;
SharedReg1071_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1071_out;
SharedReg678_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg678_out;
SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg921_out;
SharedReg162_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg162_out;
SharedReg1164_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1164_out;
SharedReg440_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg440_out;
SharedReg602_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg602_out;
SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg599_out;
SharedReg767_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg767_out;
SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg442_out;
SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg921_out;
SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg496_out;
SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg921_out;
SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg8_out;
SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg496_out;
SharedReg920_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg920_out;
SharedReg768_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg768_out;
SharedReg267_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg267_out;
SharedReg965_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg965_out;
   MUX_Add3_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1164_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg440_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg602_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg767_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg13_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg10_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg8_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg496_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg920_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg768_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg267_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg965_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg442_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg77_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg264_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1071_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg678_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg921_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg162_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_6_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_6_impl_0_out,
                 Y => Delay1No80_out);

SharedReg381_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg381_out;
SharedReg155_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg155_out;
SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg960_out;
SharedReg678_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg678_out;
SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg375_out;
SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg375_out;
SharedReg873_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg873_out;
SharedReg921_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg921_out;
SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg920_out;
SharedReg274_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg274_out;
SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg872_out;
SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg497_out;
SharedReg595_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg595_out;
SharedReg861_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg861_out;
SharedReg768_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg768_out;
SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg497_out;
SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg961_out;
SharedReg965_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg965_out;
SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg961_out;
SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg24_out;
SharedReg446_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg446_out;
SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg960_out;
SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg920_out;
SharedReg380_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg380_out;
SharedReg766_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg766_out;
   MUX_Add3_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg381_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg155_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg595_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg861_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg768_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg497_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg965_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg961_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg29_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg26_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg24_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg446_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg960_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg380_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg766_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg678_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg375_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg873_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg921_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg920_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg274_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_6_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_6_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add3_7_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add3_7_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add3_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_7_impl_out,
                 X => Delay1No82_out_to_Add3_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add3_7_impl_parent_implementedSystem_port_1_cast);

SharedReg774_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg774_out;
SharedReg280_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
SharedReg971_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg971_out;
SharedReg391_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg391_out;
SharedReg166_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg166_out;
SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg504_out;
SharedReg84_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg84_out;
SharedReg277_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg277_out;
SharedReg1084_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1084_out;
SharedReg683_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg683_out;
SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg927_out;
SharedReg172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg172_out;
SharedReg1172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1172_out;
SharedReg502_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg502_out;
SharedReg616_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg616_out;
SharedReg613_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg613_out;
SharedReg773_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg773_out;
SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg504_out;
SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg927_out;
SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg642_out;
SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg927_out;
SharedReg2_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg8_out;
SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg642_out;
SharedReg926_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg926_out;
   MUX_Add3_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg774_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg683_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1172_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg502_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg616_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg613_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg773_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg971_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg2_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg13_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg10_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg8_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg642_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg926_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg391_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg166_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg504_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg84_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg277_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1084_out_to_MUX_Add3_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_7_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_7_impl_0_out,
                 Y => Delay1No82_out);

SharedReg772_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg772_out;
SharedReg392_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg683_out;
SharedReg393_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg393_out;
SharedReg165_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg165_out;
SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg966_out;
SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg683_out;
SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg387_out;
SharedReg886_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg886_out;
SharedReg927_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg927_out;
SharedReg926_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg926_out;
SharedReg287_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg287_out;
SharedReg885_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg885_out;
SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg643_out;
SharedReg609_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg609_out;
SharedReg874_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg874_out;
SharedReg774_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg774_out;
SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg643_out;
SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg967_out;
SharedReg971_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg971_out;
SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg967_out;
SharedReg18_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg24_out;
SharedReg639_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg639_out;
SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg966_out;
   MUX_Add3_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg772_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg927_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg926_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg287_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg885_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg609_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg874_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg774_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg643_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg971_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg967_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg18_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg29_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg26_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg24_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg639_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg393_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg165_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg966_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg683_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg387_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg886_out_to_MUX_Add3_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_7_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_7_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add3_8_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add3_8_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add3_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_8_impl_out,
                 X => Delay1No84_out_to_Add3_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add3_8_impl_parent_implementedSystem_port_1_cast);

SharedReg10_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg8_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg450_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg450_out;
SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg689_out;
SharedReg691_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg691_out;
SharedReg293_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg293_out;
SharedReg978_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg978_out;
SharedReg403_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg403_out;
SharedReg176_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg452_out;
SharedReg91_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg91_out;
SharedReg290_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg290_out;
SharedReg1097_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1097_out;
SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg689_out;
SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg779_out;
SharedReg182_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg182_out;
SharedReg1180_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1180_out;
SharedReg637_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg637_out;
SharedReg630_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg630_out;
SharedReg627_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg627_out;
SharedReg727_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg727_out;
SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg452_out;
SharedReg973_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg973_out;
SharedReg505_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg505_out;
SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg779_out;
SharedReg2_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg13_out;
   MUX_Add3_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg91_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg290_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1097_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg182_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1180_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg637_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg630_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg450_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg627_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg727_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg452_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg973_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg505_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg2_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg13_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg689_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg691_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg293_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg978_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg403_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Add3_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_8_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_8_impl_0_out,
                 Y => Delay1No84_out);

SharedReg26_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg24_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg974_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg974_out;
SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg726_out;
SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg726_out;
SharedReg404_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg505_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg505_out;
SharedReg405_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg405_out;
SharedReg175_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg175_out;
SharedReg778_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg778_out;
SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg726_out;
SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg399_out;
SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg399_out;
SharedReg899_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg899_out;
SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg973_out;
SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg726_out;
SharedReg300_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg300_out;
SharedReg898_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg898_out;
SharedReg506_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg506_out;
SharedReg623_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg623_out;
SharedReg887_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg887_out;
SharedReg780_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg780_out;
SharedReg451_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg451_out;
SharedReg980_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg980_out;
SharedReg984_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg984_out;
SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg973_out;
SharedReg18_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg29_out;
   MUX_Add3_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg399_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg899_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg300_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg898_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg506_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg623_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg974_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg887_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg780_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg451_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg980_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg984_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg973_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg18_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg29_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg726_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg505_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg405_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg778_out_to_MUX_Add3_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add3_8_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_8_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No86_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg695_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg695_out;
SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1102_out;
SharedReg734_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg734_out;
SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg648_out;
SharedReg939_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg939_out;
SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg733_out;
SharedReg186_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg186_out;
SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg941_out;
SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1102_out;
SharedReg651_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg651_out;
SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg460_out;
SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg648_out;
SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1102_out;
SharedReg1105_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1105_out;
SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg648_out;
SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg648_out;
SharedReg940_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg940_out;
SharedReg306_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg306_out;
SharedReg101_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg101_out;
SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg941_out;
SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg941_out;
SharedReg411_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg411_out;
SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg733_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg186_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg651_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg460_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1105_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg15_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg940_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg306_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg101_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg941_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg411_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg733_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg11_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg695_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1102_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg734_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg648_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg939_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No86_out);

SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg732_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg940_out;
SharedReg943_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg943_out;
SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1102_out;
SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg695_out;
SharedReg1103_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1103_out;
SharedReg411_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg411_out;
SharedReg302_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg302_out;
SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1102_out;
SharedReg651_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg651_out;
SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg732_out;
SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg648_out;
SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg695_out;
SharedReg942_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg942_out;
SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1102_out;
SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg695_out;
SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg695_out;
SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1102_out;
SharedReg95_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg95_out;
SharedReg185_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg185_out;
SharedReg698_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg698_out;
SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg940_out;
SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg648_out;
SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg940_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg411_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg302_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg651_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg732_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg942_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg31_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg95_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg185_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg698_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg648_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg27_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg940_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg943_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1102_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg695_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1103_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No88_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg948_out;
SharedReg1103_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1103_out;
SharedReg702_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg14_out;
SharedReg701_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg701_out;
SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg739_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg739_out;
SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg653_out;
SharedReg946_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg946_out;
SharedReg738_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg738_out;
SharedReg199_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg199_out;
SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg948_out;
SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1106_out;
SharedReg656_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg656_out;
SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg466_out;
SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg653_out;
SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1106_out;
SharedReg1109_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1109_out;
SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg653_out;
SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg653_out;
SharedReg947_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg947_out;
SharedReg318_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg318_out;
SharedReg111_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg111_out;
SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg948_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1103_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg739_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg946_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg738_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg199_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg656_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg466_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg702_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1109_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg947_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg318_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg111_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg948_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg653_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg14_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg701_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No88_out);

SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg947_out;
SharedReg466_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg466_out;
SharedReg738_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg738_out;
SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg701_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg947_out;
SharedReg950_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg950_out;
SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1106_out;
SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg701_out;
SharedReg1107_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1107_out;
SharedReg416_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg416_out;
SharedReg314_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg314_out;
SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1106_out;
SharedReg656_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg656_out;
SharedReg737_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg737_out;
SharedReg653_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg653_out;
SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg701_out;
SharedReg949_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg949_out;
SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1106_out;
SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg701_out;
SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg701_out;
SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1106_out;
SharedReg105_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg105_out;
SharedReg198_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg198_out;
SharedReg704_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg704_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg466_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1107_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg416_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg314_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg656_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg737_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg653_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg738_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg949_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1106_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg105_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg198_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg704_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg701_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg947_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg950_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_2_impl_out,
                 X => Delay1No90_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg330_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg330_out;
SharedReg121_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg744_out;
SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg744_out;
SharedReg947_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg947_out;
SharedReg708_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg708_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg658_out;
SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg14_out;
SharedReg707_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg707_out;
SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg909_out;
SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg744_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg658_out;
SharedReg953_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg953_out;
SharedReg743_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg743_out;
SharedReg212_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg212_out;
SharedReg955_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg955_out;
SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg909_out;
SharedReg661_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg661_out;
SharedReg472_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg472_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg658_out;
SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg909_out;
SharedReg912_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg912_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg658_out;
SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg658_out;
SharedReg954_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg954_out;
   MUX_Add12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg330_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg14_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg707_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg953_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg743_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg212_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg955_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg661_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg472_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg909_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg912_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg954_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg744_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg947_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg708_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg658_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg15_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_2_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_0_out,
                 Y => Delay1No90_out);

SharedReg115_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg211_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg710_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg710_out;
SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg743_out;
SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg472_out;
SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg743_out;
SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg707_out;
SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg954_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg954_out;
SharedReg957_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg957_out;
SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg909_out;
SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg707_out;
SharedReg910_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg910_out;
SharedReg421_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg421_out;
SharedReg326_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg326_out;
SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg909_out;
SharedReg661_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg661_out;
SharedReg742_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg742_out;
SharedReg658_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg658_out;
SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg707_out;
SharedReg956_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg956_out;
SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg909_out;
SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg707_out;
SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg909_out;
   MUX_Add12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg954_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg957_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg910_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg421_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg326_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg661_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg710_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg742_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg658_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg956_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg909_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg472_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg743_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_2_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_3_impl_out,
                 X => Delay1No92_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg478_out;
SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg478_out;
SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg748_out;
SharedReg342_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg342_out;
SharedReg131_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg131_out;
SharedReg715_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg715_out;
SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg749_out;
SharedReg954_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg954_out;
SharedReg714_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg714_out;
SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg663_out;
SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg14_out;
SharedReg713_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg713_out;
SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg900_out;
SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg749_out;
SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg663_out;
SharedReg913_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg913_out;
SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg748_out;
SharedReg225_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg225_out;
SharedReg915_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg915_out;
SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg900_out;
SharedReg666_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg666_out;
SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg478_out;
SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg663_out;
SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg900_out;
Delay8No111_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast <= Delay8No111_out;
   MUX_Add12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg14_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg713_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg913_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg748_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg225_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg915_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg666_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg478_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg900_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay8No111_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg342_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg131_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg715_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg749_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg954_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg714_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg663_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_3_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_0_out,
                 Y => Delay1No92_out);

SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg663_out;
SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg663_out;
SharedReg913_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg913_out;
SharedReg125_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg224_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg666_out;
SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg748_out;
SharedReg478_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg478_out;
SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg748_out;
SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg713_out;
SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
SharedReg914_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg914_out;
SharedReg917_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg917_out;
SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg900_out;
SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg713_out;
SharedReg901_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg901_out;
SharedReg426_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg426_out;
SharedReg338_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg338_out;
SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg900_out;
SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg666_out;
SharedReg747_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg747_out;
SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg663_out;
SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg713_out;
SharedReg916_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg916_out;
SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg900_out;
   MUX_Add12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg914_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg917_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg901_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg426_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg913_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg338_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg747_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg663_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg916_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg900_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg125_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg666_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg478_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg748_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg713_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_3_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_4_impl_out,
                 X => Delay1No94_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg484_out;
SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
Delay8No112_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast <= Delay8No112_out;
SharedReg430_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg430_out;
SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg484_out;
SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg754_out;
SharedReg354_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg354_out;
SharedReg141_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg141_out;
SharedReg721_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg721_out;
SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg755_out;
SharedReg914_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg914_out;
SharedReg720_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg720_out;
SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg668_out;
SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg14_out;
SharedReg719_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg719_out;
SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg453_out;
SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg755_out;
SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg668_out;
SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg903_out;
SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg754_out;
SharedReg238_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg238_out;
SharedReg905_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg905_out;
SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg453_out;
SharedReg671_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg671_out;
SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg484_out;
   MUX_Add12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg914_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg720_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg15_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg14_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg719_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay8No112_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg668_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg903_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg238_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg905_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg453_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg671_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg430_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg484_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg754_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg354_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg141_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg721_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg755_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_4_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_0_out,
                 Y => Delay1No94_out);

SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg668_out;
SharedReg906_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg903_out;
SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg484_out;
SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg668_out;
SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg903_out;
SharedReg135_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg135_out;
SharedReg237_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg237_out;
SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg671_out;
SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg754_out;
SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg484_out;
SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg754_out;
SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg719_out;
SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg30_out;
SharedReg904_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg904_out;
SharedReg907_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg907_out;
SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg453_out;
SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg719_out;
SharedReg454_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg454_out;
SharedReg431_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg431_out;
SharedReg350_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg350_out;
SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg453_out;
SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg671_out;
SharedReg753_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg753_out;
SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg668_out;
   MUX_Add12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg31_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg30_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg904_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg907_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg719_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg454_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg431_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg350_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg453_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg753_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg484_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg668_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg135_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg237_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg671_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg754_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_4_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add12_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_5_impl_out,
                 X => Delay1No96_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast);

SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg456_out;
SharedReg676_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg676_out;
SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg435_out;
SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg435_out;
SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg456_out;
Delay8No113_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast <= Delay8No113_out;
SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg435_out;
SharedReg490_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg490_out;
SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg933_out;
SharedReg366_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg366_out;
SharedReg151_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg761_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg761_out;
SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg934_out;
SharedReg904_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg904_out;
SharedReg760_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg760_out;
SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg673_out;
SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg14_out;
SharedReg759_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg759_out;
SharedReg440_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg440_out;
SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg934_out;
SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg673_out;
SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg456_out;
SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg933_out;
SharedReg251_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg251_out;
SharedReg458_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg458_out;
   MUX_Add12_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg676_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg761_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg904_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg760_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg15_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg11_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg14_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg759_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg440_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg934_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg673_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg251_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg458_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg456_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay8No113_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg435_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg490_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg933_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg366_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_5_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_5_impl_0_out,
                 Y => Delay1No96_out);

SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg676_out;
SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg759_out;
SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg490_out;
SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg490_out;
SharedReg935_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg935_out;
SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg456_out;
SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg490_out;
SharedReg673_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg673_out;
SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg456_out;
SharedReg145_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg145_out;
SharedReg250_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg250_out;
SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg676_out;
SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg933_out;
SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg490_out;
SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg933_out;
SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg759_out;
SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg30_out;
SharedReg457_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg457_out;
SharedReg459_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg459_out;
SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg440_out;
SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg759_out;
SharedReg441_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg441_out;
SharedReg436_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg436_out;
SharedReg362_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg362_out;
SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg440_out;
   MUX_Add12_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg676_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg933_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg31_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg27_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg30_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg457_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg459_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg759_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg441_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg436_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg362_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg440_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg935_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg490_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg673_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg456_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg145_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_5_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_5_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add12_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_6_impl_out,
                 X => Delay1No98_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast);

SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg961_out;
SharedReg264_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg962_out;
SharedReg960_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg960_out;
SharedReg681_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg681_out;
SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg496_out;
SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg496_out;
SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg444_out;
SharedReg449_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg449_out;
SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg496_out;
SharedReg678_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg678_out;
SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg961_out;
SharedReg378_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg378_out;
SharedReg161_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg161_out;
SharedReg922_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg922_out;
SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg962_out;
SharedReg457_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg457_out;
SharedReg921_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg921_out;
SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg766_out;
SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg14_out;
SharedReg920_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg920_out;
SharedReg502_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg502_out;
SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg962_out;
SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg766_out;
SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg444_out;
   MUX_Add12_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg678_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg961_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg378_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg161_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg922_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg457_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg921_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg15_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg14_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg920_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg502_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg962_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg766_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg960_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg681_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg444_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg449_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg496_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_6_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_6_impl_0_out,
                 Y => Delay1No98_out);

SharedReg497_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg497_out;
SharedReg374_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg374_out;
SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg444_out;
SharedReg681_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg681_out;
SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg678_out;
SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg678_out;
SharedReg963_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg963_out;
SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg444_out;
SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg678_out;
SharedReg766_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg766_out;
SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg444_out;
SharedReg155_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg155_out;
SharedReg263_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg263_out;
SharedReg769_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg769_out;
SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg961_out;
SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg678_out;
SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg961_out;
SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg920_out;
SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg30_out;
SharedReg445_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg445_out;
SharedReg448_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg448_out;
SharedReg502_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg502_out;
SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg920_out;
SharedReg503_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg503_out;
   MUX_Add12_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg497_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg374_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg766_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg155_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg263_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg769_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg961_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg31_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg30_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg445_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg448_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg502_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg503_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg681_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg963_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg444_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg678_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_6_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_6_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add12_7_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add12_7_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add12_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_7_impl_out,
                 X => Delay1No100_out_to_Add12_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add12_7_impl_parent_implementedSystem_port_1_cast);

SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg968_out;
SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg683_out;
SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg966_out;
SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg927_out;
SharedReg277_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg277_out;
SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg928_out;
SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg966_out;
SharedReg686_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg686_out;
SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg642_out;
SharedReg637_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg637_out;
SharedReg641_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg641_out;
SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg642_out;
SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg683_out;
SharedReg967_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg967_out;
SharedReg390_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg390_out;
SharedReg171_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg171_out;
SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg928_out;
SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg968_out;
SharedReg445_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg445_out;
SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg927_out;
SharedReg772_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg772_out;
SharedReg3_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg14_out;
SharedReg926_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg926_out;
SharedReg450_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg450_out;
   MUX_Add12_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg637_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg641_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg683_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg967_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg390_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg171_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg968_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg445_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg772_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg3_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg15_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg11_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg14_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg926_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg450_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg927_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg277_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg928_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg966_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg686_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg642_out_to_MUX_Add12_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_7_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_7_impl_0_out,
                 Y => Delay1No100_out);

SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg637_out;
SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg772_out;
SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg638_out;
SharedReg503_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg503_out;
SharedReg386_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg386_out;
SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg637_out;
SharedReg645_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg645_out;
SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg926_out;
SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg683_out;
SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg683_out;
SharedReg969_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg969_out;
SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg637_out;
SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg683_out;
SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg772_out;
SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg637_out;
SharedReg165_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg165_out;
SharedReg276_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg276_out;
SharedReg775_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg775_out;
SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg967_out;
SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg683_out;
SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg967_out;
SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg926_out;
SharedReg19_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg30_out;
SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg638_out;
SharedReg640_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg640_out;
   MUX_Add12_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg969_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg772_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg165_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg276_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg775_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg967_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg19_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg31_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg27_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg30_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg638_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg640_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg503_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg386_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg637_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg645_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg926_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg683_out_to_MUX_Add12_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_7_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_7_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add12_8_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add12_8_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add12_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_8_impl_out,
                 X => Delay1No102_out_to_Add12_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add12_8_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg726_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg726_out;
SharedReg972_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg972_out;
SharedReg780_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg780_out;
SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg689_out;
SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg778_out;
SharedReg727_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg727_out;
SharedReg290_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg290_out;
SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg974_out;
SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg979_out;
SharedReg692_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg692_out;
SharedReg450_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg450_out;
SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg689_out;
SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg979_out;
SharedReg983_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg983_out;
SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg689_out;
SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg689_out;
SharedReg973_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg973_out;
SharedReg402_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg402_out;
SharedReg181_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg181_out;
SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg974_out;
SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg974_out;
SharedReg451_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg451_out;
SharedReg779_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg779_out;
SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg778_out;
SharedReg3_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg15_out;
   MUX_Add12_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg692_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg450_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg979_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg983_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg973_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg402_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg726_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg181_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg451_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg779_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg3_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg15_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg972_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg780_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg689_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg778_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg727_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg290_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg974_out_to_MUX_Add12_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_8_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_8_impl_0_out,
                 Y => Delay1No102_out);

SharedReg27_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg973_out;
SharedReg982_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg982_out;
SharedReg979_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg979_out;
SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg726_out;
SharedReg980_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg980_out;
SharedReg638_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg638_out;
SharedReg398_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg398_out;
SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg972_out;
SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg692_out;
SharedReg778_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg778_out;
SharedReg505_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg505_out;
SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg726_out;
SharedReg975_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg975_out;
SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg972_out;
SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg726_out;
SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg726_out;
SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg972_out;
SharedReg175_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg175_out;
SharedReg289_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg289_out;
SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg692_out;
SharedReg779_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg779_out;
SharedReg689_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg689_out;
SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg973_out;
SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg972_out;
SharedReg19_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg31_out;
   MUX_Add12_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg505_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg975_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg175_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg289_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg692_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg779_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg689_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg973_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg19_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg31_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg982_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg979_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg726_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg980_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg638_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg398_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg972_out_to_MUX_Add12_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Add12_8_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_8_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No104_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1194_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1197_out;
SharedReg35_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg1226_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1184_out;
SharedReg1185_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1249_out;
SharedReg514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg514_out;
SharedReg1268_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1278_out;
SharedReg1272_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1272_out;
SharedReg1200_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1201_out;
SharedReg1202_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1202_out;
SharedReg1203_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1204_out;
SharedReg1205_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1206_out;
SharedReg34_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg34_out;
SharedReg1207_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1193_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1194_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1242_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1186_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1249_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg514_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1268_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1278_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1272_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1200_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1201_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1202_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1203_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1196_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1204_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1205_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1206_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg34_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1207_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1191_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1192_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1193_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1197_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1226_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1182_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1238_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1184_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1185_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No104_out);

SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg1112_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg34_out;
SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg1225_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1225_out;
SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg34_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg783_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg783_out;
SharedReg304_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg304_out;
SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg98_out;
SharedReg188_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg188_out;
SharedReg785_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg785_out;
SharedReg1248_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1248_out;
SharedReg1115_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1115_out;
SharedReg990_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg990_out;
SharedReg991_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg991_out;
SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg186_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg33_out;
SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg95_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg33_out;
SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg186_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg33_out;
SharedReg1234_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1234_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg32_out;
SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg185_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg188_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1248_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1115_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg990_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg991_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg95_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg186_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1234_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg185_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1225_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg783_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg304_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg98_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No106_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1197_out;
SharedReg42_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg42_out;
SharedReg1226_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1184_out;
SharedReg1185_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1249_out;
SharedReg528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg528_out;
SharedReg1268_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1278_out;
SharedReg1272_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1272_out;
SharedReg1200_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1201_out;
SharedReg1202_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1202_out;
SharedReg1203_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1204_out;
SharedReg199_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg199_out;
SharedReg1206_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1235_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1192_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1238_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1184_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1185_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1186_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1249_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg528_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1268_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1278_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1272_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1200_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1193_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1201_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1202_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1203_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1204_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg199_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1206_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1209_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1235_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1194_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1242_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1197_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg42_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1226_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1182_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No106_out);

SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg1120_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg41_out;
SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg108_out;
SharedReg1225_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1225_out;
SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg41_out;
SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg39_out;
SharedReg796_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg796_out;
SharedReg316_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg316_out;
SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg108_out;
SharedReg201_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg201_out;
SharedReg798_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg798_out;
SharedReg1248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1248_out;
SharedReg1123_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1123_out;
SharedReg1003_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1003_out;
SharedReg1004_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1004_out;
SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg105_out;
SharedReg199_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg199_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg40_out;
SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg105_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg40_out;
SharedReg1232_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1232_out;
SharedReg107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg107_out;
SharedReg113_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg113_out;
SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg39_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg796_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg316_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg201_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg798_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1123_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1003_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1004_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg199_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg105_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1232_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg113_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg198_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg108_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1225_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg41_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No108_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1206_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1197_out;
SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg49_out;
SharedReg1226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1184_out;
SharedReg1185_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1249_out;
SharedReg542_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg542_out;
SharedReg1268_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1278_out;
SharedReg1272_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1272_out;
SharedReg1200_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1229_out;
SharedReg115_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg115_out;
SharedReg1231_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1205_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1206_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1209_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg49_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1226_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1182_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1238_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1184_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1185_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1186_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1249_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg542_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1268_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1235_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1278_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1272_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1200_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1201_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1229_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg115_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1231_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1205_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1191_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1192_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1193_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1194_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1242_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1196_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1197_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No108_out);

SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg123_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg46_out;
SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg46_out;
SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg211_out;
SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg211_out;
SharedReg1128_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1128_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg48_out;
SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg118_out;
SharedReg1225_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1225_out;
SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg48_out;
SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg46_out;
SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg809_out;
SharedReg328_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg328_out;
SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg118_out;
SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg214_out;
SharedReg811_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg811_out;
SharedReg1248_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1248_out;
SharedReg1131_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1131_out;
SharedReg1016_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1016_out;
SharedReg1017_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1017_out;
SharedReg115_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg115_out;
SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg212_out;
SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg47_out;
SharedReg1230_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1230_out;
SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg47_out;
SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg47_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1225_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg328_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg811_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1248_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1131_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1016_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1017_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg115_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1230_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg47_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg46_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1128_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg48_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No110_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg125_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg1231_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1197_out;
SharedReg56_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg56_out;
SharedReg1226_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1184_out;
SharedReg1185_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1249_out;
SharedReg556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg556_out;
SharedReg1268_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1278_out;
SharedReg1252_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1227_out;
SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg225_out;
SharedReg53_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg53_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1231_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1242_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1196_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1197_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg56_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1226_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1184_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1185_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1186_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1205_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1249_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg556_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1268_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1278_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1252_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1227_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg225_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg53_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1206_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1209_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1235_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1191_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1192_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1193_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1194_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No110_out);

SharedReg1230_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1230_out;
SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg54_out;
SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg127_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg133_out;
SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg53_out;
SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg53_out;
SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg53_out;
SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg224_out;
SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg224_out;
SharedReg1136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1136_out;
SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg55_out;
SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg128_out;
SharedReg1225_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1225_out;
SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg55_out;
SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg53_out;
SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg822_out;
SharedReg340_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg340_out;
SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg128_out;
SharedReg227_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg227_out;
SharedReg824_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg824_out;
SharedReg1248_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1248_out;
SharedReg1139_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1139_out;
SharedReg1029_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1029_out;
SharedReg1033_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1033_out;
SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg125_out;
SharedReg1228_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1229_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1230_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1136_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1225_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg55_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg340_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg128_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg227_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg54_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg824_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1248_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1139_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1029_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1033_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1228_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1229_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg127_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg53_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg224_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No112_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1227_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1227_out;
SharedReg238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg60_out;
SharedReg135_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg135_out;
SharedReg1231_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1197_out;
SharedReg63_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg63_out;
SharedReg1226_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1184_out;
SharedReg1185_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1247_out;
SharedReg1147_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1147_out;
SharedReg1190_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1252_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1227_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1192_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1193_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1242_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1197_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg63_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1226_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1182_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1238_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1184_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1185_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1186_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1249_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1247_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1147_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1190_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1252_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg135_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1231_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1205_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1206_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1209_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1235_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No112_out);

SharedReg135_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg1228_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1229_out;
SharedReg1230_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1230_out;
SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg61_out;
SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg61_out;
SharedReg137_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg137_out;
SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg143_out;
SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg60_out;
SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg60_out;
SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg237_out;
SharedReg1144_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1144_out;
SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg62_out;
SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg138_out;
SharedReg1225_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1225_out;
SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg60_out;
SharedReg835_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg835_out;
SharedReg352_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg352_out;
SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg138_out;
SharedReg240_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg240_out;
SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg837_out;
SharedReg571_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg571_out;
SharedReg1270_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1270_out;
SharedReg241_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg241_out;
SharedReg1047_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1047_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1228_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg237_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1144_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1225_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg835_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1229_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg352_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg138_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg240_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg571_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1270_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg241_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1047_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1230_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg61_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg137_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg60_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product4_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_5_impl_out,
                 X => Delay1No114_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1155_out;
SharedReg1190_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1227_out;
SharedReg251_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg251_out;
SharedReg67_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg145_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg145_out;
SharedReg1231_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1197_out;
SharedReg70_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg70_out;
SharedReg1226_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1226_out;
SharedReg1182_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1184_out;
SharedReg148_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg148_out;
SharedReg1267_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1247_out;
   MUX_Product4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1190_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1209_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1235_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1191_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1192_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1193_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1194_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1242_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1196_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1197_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg70_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1252_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1226_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1182_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1238_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1184_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg148_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1267_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1249_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1247_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1227_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg251_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg145_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1231_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1205_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1206_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_5_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_0_out,
                 Y => Delay1No114_out);

SharedReg1270_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1270_out;
SharedReg254_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg254_out;
SharedReg1060_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1060_out;
SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg1228_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1229_out;
SharedReg1230_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1230_out;
SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg68_out;
SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg147_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg147_out;
SharedReg153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg153_out;
SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg67_out;
SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg67_out;
SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg67_out;
SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg250_out;
SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg250_out;
SharedReg1152_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1152_out;
SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg69_out;
SharedReg148_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg148_out;
SharedReg1225_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1225_out;
SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg69_out;
SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg67_out;
SharedReg848_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg848_out;
SharedReg364_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg364_out;
SharedReg1213_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1213_out;
SharedReg1052_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1052_out;
SharedReg851_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg851_out;
SharedReg584_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg584_out;
   MUX_Product4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1270_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg250_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1152_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg148_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1225_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1060_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg69_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg67_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg848_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg364_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1213_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1052_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg851_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg584_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1228_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1229_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1230_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg147_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_5_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product4_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_6_impl_out,
                 X => Delay1No116_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1247_out;
SharedReg1268_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1278_out;
SharedReg1252_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1229_out;
SharedReg1203_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1204_out;
SharedReg264_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg264_out;
SharedReg1206_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1206_out;
SharedReg76_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg76_out;
SharedReg1207_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1207_out;
SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1150_out;
SharedReg1153_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1153_out;
SharedReg1275_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1259_out;
SharedReg1152_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1152_out;
SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1150_out;
SharedReg1183_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1288_out;
SharedReg1182_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1184_out;
SharedReg158_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg158_out;
   MUX_Product4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1249_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1204_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg264_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1206_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg76_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1207_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1153_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1275_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1281_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1259_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1247_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1152_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1183_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1288_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1182_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1238_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1184_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg158_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1268_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1278_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1252_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1200_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1201_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1229_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1203_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_6_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_0_out,
                 Y => Delay1No116_out);

SharedReg266_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg863_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg863_out;
SharedReg599_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg599_out;
SharedReg1163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1163_out;
SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1068_out;
SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1072_out;
SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg264_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg264_out;
SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg75_out;
SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg155_out;
SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg75_out;
SharedReg1232_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1232_out;
SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg75_out;
SharedReg1234_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1234_out;
SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg74_out;
SharedReg1245_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1280_out;
SharedReg1154_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1154_out;
SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1152_out;
SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1152_out;
SharedReg1260_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1287_out;
SharedReg250_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg250_out;
SharedReg1052_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1052_out;
SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg74_out;
SharedReg861_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg861_out;
SharedReg376_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg376_out;
SharedReg1213_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1213_out;
   MUX_Product4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg863_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1232_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1234_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1245_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1280_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1154_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1152_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg599_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1260_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1287_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg250_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1052_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg74_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg861_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg376_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1213_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1072_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg264_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg75_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg155_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_6_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product4_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_7_impl_out,
                 X => Delay1No118_out_to_Product4_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product4_7_impl_parent_implementedSystem_port_1_cast);

SharedReg377_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg377_out;
SharedReg1187_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1187_out;
SharedReg1185_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1185_out;
SharedReg1189_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1218_out;
SharedReg612_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg612_out;
SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1263_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1272_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1272_out;
SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg863_out;
SharedReg1160_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1160_out;
SharedReg1202_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1202_out;
SharedReg1161_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1161_out;
SharedReg1165_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1165_out;
SharedReg1205_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1205_out;
SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1063_out;
SharedReg1279_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1245_out;
SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg863_out;
SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg863_out;
SharedReg1276_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1251_out;
SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1158_out;
SharedReg1183_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1288_out;
SharedReg1182_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1182_out;
   MUX_Product4_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg377_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1187_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1160_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1202_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1161_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1165_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1205_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1063_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1279_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1244_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1245_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1185_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1276_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1250_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1251_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1183_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1288_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1182_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1189_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1218_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg612_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1272_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg863_out_to_MUX_Product4_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_7_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_7_impl_0_out,
                 Y => Delay1No118_out);

SharedReg1214_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1214_out;
SharedReg600_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg600_out;
SharedReg168_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg379_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg79_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg79_out;
SharedReg1248_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1248_out;
SharedReg1262_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1262_out;
SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1064_out;
SharedReg1082_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1082_out;
SharedReg1265_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1231_out;
SharedReg82_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg82_out;
SharedReg1233_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1237_out;
SharedReg277_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg277_out;
SharedReg1219_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1219_out;
SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1063_out;
SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1063_out;
SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1063_out;
SharedReg1280_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1223_out;
SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1160_out;
SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1160_out;
SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1160_out;
SharedReg1287_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1287_out;
SharedReg263_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg263_out;
SharedReg1065_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1065_out;
SharedReg81_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg81_out;
   MUX_Product4_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1214_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg600_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1231_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg82_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1233_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1237_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg277_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1219_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1063_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1280_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1223_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1160_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1287_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg263_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1065_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg81_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg379_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg79_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1248_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1262_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1064_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1082_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1265_out_to_MUX_Product4_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_7_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_7_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product4_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_8_impl_out,
                 X => Delay1No120_out_to_Product4_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product4_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1197_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1197_out;
SharedReg91_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg1199_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1199_out;
SharedReg1182_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1182_out;
SharedReg1238_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1238_out;
SharedReg1212_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1212_out;
SharedReg1185_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1249_out;
SharedReg626_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg626_out;
SharedReg1268_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1268_out;
SharedReg1190_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1190_out;
SharedReg1272_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1272_out;
SharedReg1200_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1200_out;
SharedReg290_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg290_out;
SharedReg1202_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1202_out;
SharedReg1203_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1203_out;
SharedReg1231_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1206_out;
SharedReg90_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg90_out;
SharedReg1166_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1166_out;
SharedReg1169_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1169_out;
SharedReg1275_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1275_out;
SharedReg1193_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1242_out;
SharedReg1223_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1223_out;
   MUX_Product4_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1197_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1268_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1190_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1272_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1200_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg290_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1202_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1203_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1231_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1205_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1206_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1199_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg90_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1166_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1169_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1275_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1193_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1194_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1242_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1223_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1182_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1238_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1212_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1185_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1186_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1249_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg626_out_to_MUX_Product4_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_8_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_8_impl_0_out,
                 Y => Delay1No120_out);

SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg1225_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1225_out;
SharedReg895_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg895_out;
SharedReg88_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg88_out;
SharedReg887_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg887_out;
SharedReg291_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg291_out;
SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg292_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg292_out;
SharedReg890_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg890_out;
SharedReg1248_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1248_out;
SharedReg1179_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1179_out;
SharedReg293_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg293_out;
SharedReg1095_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1095_out;
SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg175_out;
SharedReg1228_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1228_out;
SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg89_out;
SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg175_out;
SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg89_out;
SharedReg290_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg290_out;
SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg89_out;
SharedReg1234_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1234_out;
SharedReg1245_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1280_out;
SharedReg1170_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1170_out;
SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg289_out;
SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg289_out;
SharedReg1176_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1176_out;
SharedReg90_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg90_out;
   MUX_Product4_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1225_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1179_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg293_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1095_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1228_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg175_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg290_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg89_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg895_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1234_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1245_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1280_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1170_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg289_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1176_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg90_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg88_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg887_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg291_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg292_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg890_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1248_out_to_MUX_Product4_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product4_8_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_8_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product11_5_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product11_5_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product11_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_5_impl_out,
                 X => Delay1No122_out_to_Product11_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product11_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1268_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1278_out;
SharedReg1252_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1229_out;
SharedReg1203_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1204_out;
SharedReg251_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg251_out;
SharedReg1206_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1206_out;
SharedReg69_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg69_out;
SharedReg1207_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1207_out;
SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1142_out;
SharedReg1145_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1145_out;
SharedReg1275_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1259_out;
SharedReg1144_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1144_out;
SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1142_out;
SharedReg1183_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1288_out;
SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1185_out;
SharedReg353_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg353_out;
SharedReg1187_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1187_out;
SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1185_out;
SharedReg1186_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1247_out;
   MUX_Product11_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1268_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1278_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg69_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1207_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1145_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1275_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1281_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1259_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1144_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1142_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1183_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1252_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1288_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg353_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1187_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1185_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1186_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1249_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1247_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1200_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1201_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1229_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1203_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1204_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg251_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1206_out_to_MUX_Product11_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_5_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_5_impl_0_out,
                 Y => Delay1No122_out);

SharedReg1155_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1155_out;
SharedReg1055_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1055_out;
SharedReg1059_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1059_out;
SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg145_out;
SharedReg251_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg251_out;
SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg68_out;
SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg145_out;
SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg68_out;
SharedReg1232_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1232_out;
SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg68_out;
SharedReg1234_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1234_out;
SharedReg67_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg67_out;
SharedReg1245_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1280_out;
SharedReg1146_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1146_out;
SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1144_out;
SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1144_out;
SharedReg1260_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1287_out;
SharedReg237_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg237_out;
SharedReg1039_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1039_out;
SharedReg838_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg838_out;
SharedReg1214_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1214_out;
SharedReg572_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg572_out;
SharedReg148_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg148_out;
SharedReg253_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg253_out;
SharedReg850_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg850_out;
SharedReg585_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg585_out;
   MUX_Product11_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1155_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1055_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1234_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg67_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1245_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1280_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1146_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1144_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1260_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1287_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg237_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1059_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1039_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg838_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1214_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg572_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg148_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg253_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg850_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg585_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg251_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg145_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1232_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg68_out_to_MUX_Product11_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_5_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_5_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product11_6_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product11_6_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product11_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_6_impl_out,
                 X => Delay1No124_out_to_Product11_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product11_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1189_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1218_out;
SharedReg598_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg598_out;
SharedReg1150_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1150_out;
SharedReg1263_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1263_out;
SharedReg1272_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1272_out;
SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg850_out;
SharedReg1152_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1152_out;
SharedReg1202_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1202_out;
SharedReg1153_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1153_out;
SharedReg1157_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1157_out;
SharedReg1205_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1205_out;
SharedReg1050_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1050_out;
SharedReg1279_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1245_out;
SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg850_out;
SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg850_out;
SharedReg1276_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1286_out;
SharedReg145_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg145_out;
SharedReg1212_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1212_out;
SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1185_out;
SharedReg365_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg365_out;
SharedReg1187_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1187_out;
SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1185_out;
   MUX_Product11_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1189_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1218_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1157_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1205_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1050_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1279_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1244_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1245_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1276_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1250_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg598_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1251_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1286_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg145_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1212_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg365_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1187_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1185_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1150_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1263_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1272_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg850_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1152_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1202_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1153_out_to_MUX_Product11_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_6_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_6_impl_0_out,
                 Y => Delay1No124_out);

SharedReg367_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg72_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg1248_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1248_out;
SharedReg1262_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1262_out;
SharedReg1051_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1051_out;
SharedReg1069_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1069_out;
SharedReg1265_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1231_out;
SharedReg75_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg75_out;
SharedReg1233_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1237_out;
SharedReg264_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg264_out;
SharedReg1219_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1219_out;
SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1050_out;
SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1050_out;
SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1050_out;
SharedReg1280_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1223_out;
SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1152_out;
SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1152_out;
SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1152_out;
SharedReg1150_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1150_out;
SharedReg1211_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1211_out;
SharedReg68_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg68_out;
SharedReg851_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg851_out;
SharedReg1214_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1214_out;
SharedReg586_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg586_out;
SharedReg158_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg158_out;
   MUX_Product11_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1237_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg264_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1219_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1050_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1280_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1223_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1248_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1152_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1150_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1211_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg68_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg851_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1214_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg586_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg158_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1262_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1051_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1069_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1265_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1231_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg75_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1233_out_to_MUX_Product11_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product11_6_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_6_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1194_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1194_out;
SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg1223_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1223_out;
SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg1198_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1212_out;
SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg98_out;
SharedReg1267_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1247_out;
SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1115_out;
SharedReg1190_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1227_out;
SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg186_out;
SharedReg1229_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1229_out;
SharedReg95_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg95_out;
SharedReg1231_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1231_out;
SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg186_out;
SharedReg1206_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1193_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1194_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1267_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1249_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1247_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1190_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1252_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1227_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1229_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg95_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1223_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1231_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg186_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1206_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1209_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1235_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1191_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1192_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1193_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1198_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1199_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1210_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1271_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1212_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No126_out);

SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg1246_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1246_out;
SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg34_out;
SharedReg1224_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1224_out;
SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg791_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg985_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg985_out;
SharedReg187_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg187_out;
SharedReg1213_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1213_out;
SharedReg987_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg987_out;
SharedReg786_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg786_out;
SharedReg515_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg515_out;
SharedReg1270_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1270_out;
SharedReg189_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg189_out;
SharedReg994_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg994_out;
SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg95_out;
SharedReg1228_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1228_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg33_out;
SharedReg1230_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1230_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg33_out;
SharedReg1232_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1232_out;
SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg97_out;
SharedReg103_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg103_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg32_out;
SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg95_out;
SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg302_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1246_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg987_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg786_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg515_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1270_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg189_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg994_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1228_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1230_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1232_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg103_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg302_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1224_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg985_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg187_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1213_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No128_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1194_out;
SharedReg1120_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg1223_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1223_out;
SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg108_out;
SharedReg1198_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1212_out;
SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg108_out;
SharedReg1267_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1247_out;
SharedReg1123_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1123_out;
SharedReg1190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1227_out;
SharedReg199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg199_out;
SharedReg1229_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1229_out;
SharedReg105_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg105_out;
SharedReg1231_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1233_out;
SharedReg113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg113_out;
SharedReg1207_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1207_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1192_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1271_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1212_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1267_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1249_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1247_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1123_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1252_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1227_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1229_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg105_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1231_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1205_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1233_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1207_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1223_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1198_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1199_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1210_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No128_out);

SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg314_out;
SharedReg1246_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1246_out;
SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg41_out;
SharedReg1224_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1224_out;
SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg107_out;
SharedReg804_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg804_out;
SharedReg39_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg39_out;
SharedReg998_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg998_out;
SharedReg200_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg200_out;
SharedReg1213_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1213_out;
SharedReg1000_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1000_out;
SharedReg799_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg799_out;
SharedReg529_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg529_out;
SharedReg1270_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1270_out;
SharedReg202_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg202_out;
SharedReg1007_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1007_out;
SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg105_out;
SharedReg1228_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1228_out;
SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg40_out;
SharedReg1230_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1230_out;
SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg40_out;
SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg40_out;
SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg107_out;
SharedReg1237_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1237_out;
SharedReg1119_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1119_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg998_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg200_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1213_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1000_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg799_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg529_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1270_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg202_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1007_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg105_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1228_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1230_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg40_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1237_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1119_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg314_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1246_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg41_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1224_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg107_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg804_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg39_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No130_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1233_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1233_out;
SharedReg123_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg1207_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1194_out;
SharedReg1128_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1128_out;
SharedReg1223_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1223_out;
SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg118_out;
SharedReg1198_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1212_out;
SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg118_out;
SharedReg1267_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1247_out;
SharedReg1131_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1131_out;
SharedReg1190_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1227_out;
SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg212_out;
SharedReg46_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg46_out;
SharedReg1203_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1232_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1233_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1198_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1199_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1271_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1267_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1249_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1247_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1131_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1207_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1190_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1252_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1227_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg46_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1203_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1204_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1232_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1191_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1192_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1193_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1194_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1128_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1223_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No130_out);

SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg1237_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1237_out;
SharedReg1127_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1127_out;
SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg115_out;
SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg326_out;
SharedReg1246_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1246_out;
SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg48_out;
SharedReg1224_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1224_out;
SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg117_out;
SharedReg817_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg817_out;
SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg46_out;
SharedReg1011_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1011_out;
SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg213_out;
SharedReg1213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1213_out;
SharedReg1013_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1013_out;
SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg812_out;
SharedReg543_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg543_out;
SharedReg1270_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1270_out;
SharedReg215_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg215_out;
SharedReg1020_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1020_out;
SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg115_out;
SharedReg1228_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1229_out;
SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg47_out;
SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg212_out;
SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg47_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1237_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg117_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg817_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1011_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1013_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg543_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1270_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1127_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg215_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1020_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1228_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1229_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg47_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg115_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1246_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg48_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1224_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No132_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1203_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1233_out;
SharedReg133_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg133_out;
SharedReg1207_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1194_out;
SharedReg1136_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1136_out;
SharedReg1223_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1223_out;
SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg128_out;
SharedReg1198_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1212_out;
SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg128_out;
SharedReg1267_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1247_out;
SharedReg1139_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1139_out;
SharedReg1190_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1255_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1203_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1204_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1136_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1223_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1198_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1199_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1210_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1271_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1212_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg128_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1267_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1249_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1247_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1139_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1190_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1252_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1200_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1254_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1255_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg133_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1207_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1191_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1192_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1193_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1194_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No132_out);

SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg225_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg225_out;
SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg1237_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1237_out;
SharedReg1135_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1135_out;
SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg125_out;
SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg125_out;
SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg338_out;
SharedReg1246_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1246_out;
SharedReg55_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg55_out;
SharedReg1224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1224_out;
SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
SharedReg830_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg830_out;
SharedReg53_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg53_out;
SharedReg1024_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1024_out;
SharedReg226_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg226_out;
SharedReg1213_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1213_out;
SharedReg1026_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1026_out;
SharedReg825_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg825_out;
SharedReg557_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg557_out;
SharedReg1270_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1270_out;
SharedReg228_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg228_out;
SharedReg1034_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1034_out;
SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg338_out;
SharedReg554_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg554_out;
SharedReg1025_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1025_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg225_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1246_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg55_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1224_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg830_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg53_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1024_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg226_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1213_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1026_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg54_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg825_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg557_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1270_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg228_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1034_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg554_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1025_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1237_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1135_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg125_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg338_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product21_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_4_impl_out,
                 X => Delay1No134_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1200_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1255_out;
SharedReg1203_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1233_out;
SharedReg143_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg143_out;
SharedReg1207_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1194_out;
SharedReg1144_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1144_out;
SharedReg1223_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1223_out;
SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg138_out;
SharedReg1198_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1212_out;
SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg138_out;
SharedReg1267_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1261_out;
   MUX_Product21_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1200_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1254_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1192_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1193_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1194_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1144_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1223_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1198_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1199_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1210_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1271_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1255_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1212_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg138_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1267_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1249_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1247_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1189_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1218_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1261_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1203_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1204_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1232_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1233_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg143_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1207_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1191_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_4_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_0_out,
                 Y => Delay1No134_out);

SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg568_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg1038_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1038_out;
SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg61_out;
SharedReg238_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg238_out;
SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg61_out;
SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg137_out;
SharedReg1237_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1237_out;
SharedReg1143_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1143_out;
SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg135_out;
SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg135_out;
SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg350_out;
SharedReg1246_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1246_out;
SharedReg62_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg62_out;
SharedReg1224_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1224_out;
SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg137_out;
SharedReg843_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg843_out;
SharedReg60_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg60_out;
SharedReg1037_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1037_out;
SharedReg239_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg239_out;
SharedReg1213_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1213_out;
SharedReg1039_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1039_out;
SharedReg838_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg838_out;
SharedReg570_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg570_out;
SharedReg139_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg139_out;
SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg241_out;
SharedReg1046_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1046_out;
   MUX_Product21_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg350_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1246_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg62_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1224_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg843_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg60_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1037_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1038_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg239_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1213_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1039_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg838_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg570_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg139_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1046_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg238_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg137_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1237_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1143_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg135_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_4_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product21_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_5_impl_out,
                 X => Delay1No136_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1189_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1261_out;
SharedReg1200_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1255_out;
SharedReg1203_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1233_out;
SharedReg153_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg153_out;
SharedReg1207_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1194_out;
SharedReg1152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1152_out;
SharedReg1223_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1223_out;
SharedReg148_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg148_out;
SharedReg1198_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1212_out;
SharedReg1239_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1258_out;
SharedReg1248_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1248_out;
   MUX_Product21_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1189_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1218_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg153_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1207_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1191_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1192_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1193_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1194_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1223_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg148_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1198_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1261_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1199_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1210_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1271_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1212_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1239_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1269_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1258_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1248_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1200_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1254_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1255_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1203_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1204_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1232_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1233_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_5_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_5_impl_0_out,
                 Y => Delay1No136_out);

SharedReg149_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg254_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg254_out;
SharedReg1059_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1059_out;
SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg362_out;
SharedReg582_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg582_out;
SharedReg1051_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1051_out;
SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg68_out;
SharedReg251_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg251_out;
SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg147_out;
SharedReg1237_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1237_out;
SharedReg1151_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1151_out;
SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg145_out;
SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg145_out;
SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg362_out;
SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg362_out;
SharedReg1246_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1246_out;
SharedReg69_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg69_out;
SharedReg1224_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1224_out;
SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg147_out;
SharedReg856_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg856_out;
SharedReg67_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg67_out;
SharedReg1050_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1050_out;
SharedReg252_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg252_out;
SharedReg583_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg583_out;
SharedReg1052_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1052_out;
SharedReg850_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg850_out;
SharedReg585_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg585_out;
   MUX_Product21_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1237_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1151_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1246_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg69_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1224_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1059_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg856_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg67_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1050_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg252_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg583_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1052_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg850_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg585_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg362_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg582_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1051_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg251_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg147_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_5_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_5_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product21_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_6_impl_out,
                 X => Delay1No138_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1267_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1247_out;
SharedReg1163_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1163_out;
SharedReg1190_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1227_out;
SharedReg264_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg264_out;
SharedReg74_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg74_out;
SharedReg155_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg155_out;
SharedReg1231_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1197_out;
SharedReg77_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg77_out;
SharedReg1226_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1212_out;
SharedReg1239_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1239_out;
   MUX_Product21_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1267_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1249_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1231_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1205_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1206_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1209_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1235_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1191_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1192_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1193_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1194_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1242_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1247_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1196_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1197_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg77_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1226_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1210_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1271_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1212_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1239_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1163_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1190_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1252_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1227_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg264_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg74_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg155_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_6_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_6_impl_0_out,
                 Y => Delay1No138_out);

SharedReg1065_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1065_out;
SharedReg864_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg864_out;
SharedReg598_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg598_out;
SharedReg1270_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1270_out;
SharedReg267_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg267_out;
SharedReg1073_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1073_out;
SharedReg155_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg155_out;
SharedReg1228_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1229_out;
SharedReg1230_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1230_out;
SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg75_out;
SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg75_out;
SharedReg157_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg157_out;
SharedReg163_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg163_out;
SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg74_out;
SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg74_out;
SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg74_out;
SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg263_out;
SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg263_out;
SharedReg1160_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1160_out;
SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg76_out;
SharedReg158_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg158_out;
SharedReg1225_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1225_out;
SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg76_out;
SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg74_out;
SharedReg1063_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1063_out;
SharedReg265_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg265_out;
SharedReg597_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg597_out;
   MUX_Product21_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1065_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg864_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg75_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg157_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg163_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg263_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1160_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg598_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg158_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1225_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg76_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg74_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1063_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg265_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg597_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1270_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1073_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg155_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1228_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1229_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1230_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_6_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_6_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product21_7_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product21_7_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product21_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_7_impl_out,
                 X => Delay1No140_out_to_Product21_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product21_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1238_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1238_out;
SharedReg1184_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1184_out;
SharedReg168_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg1186_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1186_out;
SharedReg1249_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1247_out;
SharedReg1268_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1278_out;
SharedReg1252_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1229_out;
SharedReg1203_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1204_out;
SharedReg277_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg277_out;
SharedReg1206_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1206_out;
SharedReg83_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg83_out;
SharedReg1207_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1207_out;
SharedReg1158_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1158_out;
SharedReg1161_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1161_out;
SharedReg1275_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1259_out;
SharedReg1160_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1160_out;
SharedReg1197_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1197_out;
SharedReg84_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg84_out;
SharedReg1226_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1210_out;
   MUX_Product21_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1238_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1184_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1201_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1229_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1203_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1204_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg277_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1206_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg83_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1207_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1158_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1161_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1275_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1281_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1259_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1160_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1197_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg84_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1226_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1210_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1186_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1249_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1247_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1268_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1278_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1252_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1200_out_to_MUX_Product21_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_7_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_7_impl_0_out,
                 Y => Delay1No140_out);

SharedReg874_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg874_out;
SharedReg388_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg1213_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1213_out;
SharedReg279_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg279_out;
SharedReg876_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg876_out;
SharedReg613_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg613_out;
SharedReg1171_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1171_out;
SharedReg1081_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1081_out;
SharedReg1085_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1085_out;
SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg165_out;
SharedReg277_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg277_out;
SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg82_out;
SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg82_out;
SharedReg1232_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1232_out;
SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg82_out;
SharedReg1234_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1234_out;
SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg81_out;
SharedReg1245_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1280_out;
SharedReg1162_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1162_out;
SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1160_out;
SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1160_out;
SharedReg1260_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1260_out;
SharedReg168_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg168_out;
SharedReg1225_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1225_out;
SharedReg83_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg83_out;
SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg81_out;
   MUX_Product21_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg874_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg277_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1232_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg82_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1234_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1245_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1280_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1213_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1162_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1160_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1260_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg168_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1225_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg83_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg81_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg279_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg876_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg613_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1171_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1081_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1085_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg165_out_to_MUX_Product21_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_7_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_7_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product21_8_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product21_8_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product21_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_8_impl_out,
                 X => Delay1No142_out_to_Product21_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product21_8_impl_parent_implementedSystem_port_1_cast);

SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg1198_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1210_out;
SharedReg1271_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1271_out;
SharedReg400_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg1267_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1267_out;
SharedReg1258_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1258_out;
SharedReg1247_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1247_out;
SharedReg1179_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1179_out;
SharedReg1218_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1218_out;
SharedReg1252_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1227_out;
SharedReg1254_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1254_out;
SharedReg1229_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1229_out;
SharedReg175_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg175_out;
SharedReg1204_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1204_out;
SharedReg290_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg290_out;
SharedReg1206_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1194_out;
SharedReg1176_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1176_out;
SharedReg1196_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1196_out;
   MUX_Product21_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1198_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1179_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1218_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1252_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1227_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1254_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1229_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg175_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1204_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg290_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1206_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1226_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1209_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1207_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1191_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1192_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1193_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1194_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1176_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1196_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1210_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1271_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1267_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1258_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1247_out_to_MUX_Product21_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_8_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_8_impl_0_out,
                 Y => Delay1No142_out);

SharedReg1224_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1224_out;
SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg177_out;
SharedReg895_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg895_out;
SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg88_out;
SharedReg1089_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1089_out;
SharedReg1212_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1212_out;
SharedReg1213_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1213_out;
SharedReg1091_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1091_out;
SharedReg889_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg889_out;
SharedReg627_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg627_out;
SharedReg1270_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1270_out;
SharedReg293_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg293_out;
SharedReg1098_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1098_out;
SharedReg175_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg175_out;
SharedReg624_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg624_out;
SharedReg89_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg89_out;
SharedReg1230_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1230_out;
SharedReg290_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg290_out;
SharedReg1232_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1232_out;
SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg177_out;
SharedReg183_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg183_out;
SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg88_out;
SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg88_out;
SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg88_out;
SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg398_out;
SharedReg1246_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1246_out;
SharedReg625_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg625_out;
   MUX_Product21_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1224_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1270_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg293_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1098_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg175_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg624_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg89_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1230_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg290_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1232_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg177_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg895_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg183_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg398_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1246_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg625_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg88_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1089_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1212_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1213_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1091_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg889_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg627_out_to_MUX_Product21_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product21_8_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_8_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No144_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg410_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg411_out;
Delay6No90_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= Delay6No90_out;
SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg411_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg460_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg460_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg732_out;
SharedReg784_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg784_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg732_out;
SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg413_out;
SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg410_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg460_out;
SharedReg463_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg463_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg460_out;
SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg410_out;
SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg311_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg732_out;
SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg412_out;
SharedReg516_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg516_out;
SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg412_out;
SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg411_out;
SharedReg649_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg649_out;
SharedReg461_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg461_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg784_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg463_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg410_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg732_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg516_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg412_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg649_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg461_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay6No90_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg411_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg460_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No144_out);

SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg696_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg696_out;
SharedReg700_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg700_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg460_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg732_out;
SharedReg945_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg945_out;
SharedReg1102_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1102_out;
SharedReg783_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg783_out;
SharedReg940_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg940_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg460_out;
SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg650_out;
SharedReg695_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg695_out;
SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg410_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg460_out;
SharedReg942_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg942_out;
Delay8No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast <= Delay8No36_out;
SharedReg312_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg312_out;
SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg733_out;
SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg461_out;
SharedReg511_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg511_out;
SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg650_out;
SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg462_out;
SharedReg697_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg697_out;
SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg462_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1102_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg783_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg940_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg695_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg942_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay8No36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg312_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg461_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg511_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg650_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg697_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg696_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg700_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg945_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No146_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg416_out;
SharedReg467_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg467_out;
SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg416_out;
SharedReg1102_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1102_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg416_out;
Delay6No91_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= Delay6No91_out;
SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg416_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg466_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg466_out;
SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg737_out;
SharedReg797_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg797_out;
SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg737_out;
SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg418_out;
SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg415_out;
SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg415_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg466_out;
SharedReg469_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg469_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg466_out;
SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg415_out;
SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg323_out;
SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg737_out;
SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg417_out;
SharedReg530_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg530_out;
SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg417_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg467_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg797_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg469_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg466_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg415_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg737_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg530_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg417_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1102_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg416_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay6No91_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No146_out);

SharedReg468_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg468_out;
SharedReg703_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg703_out;
SharedReg417_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg417_out;
SharedReg1103_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1103_out;
SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg702_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg702_out;
SharedReg706_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg706_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg466_out;
SharedReg737_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg737_out;
SharedReg952_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg952_out;
SharedReg1106_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1106_out;
SharedReg796_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg796_out;
SharedReg947_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg947_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg466_out;
SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg655_out;
SharedReg701_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg701_out;
SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg415_out;
SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg466_out;
SharedReg949_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg949_out;
Delay8No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast <= Delay8No37_out;
SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg324_out;
SharedReg738_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg738_out;
SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg467_out;
SharedReg525_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg525_out;
SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg655_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg468_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg703_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg737_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg952_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1106_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg796_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg947_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg701_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg417_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg466_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg949_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay8No37_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg738_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg525_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg655_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1103_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg702_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg706_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No148_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg422_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg544_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg544_out;
SharedReg1108_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1108_out;
SharedReg1107_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg421_out;
SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg421_out;
SharedReg1106_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg7_out;
SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg421_out;
Delay6No92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= Delay6No92_out;
SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg421_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg472_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg472_out;
SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg742_out;
SharedReg810_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg810_out;
SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg742_out;
SharedReg423_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg423_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg420_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg420_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg472_out;
SharedReg475_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg475_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg472_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg420_out;
SharedReg335_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg335_out;
SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg742_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg544_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay6No92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg810_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg423_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1108_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg475_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg335_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg742_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No148_out);

SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg473_out;
SharedReg539_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg539_out;
SharedReg474_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg474_out;
SharedReg422_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg422_out;
SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg660_out;
SharedReg1108_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1108_out;
SharedReg1107_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1107_out;
SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg23_out;
SharedReg708_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg708_out;
SharedReg712_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg712_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg472_out;
SharedReg742_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg742_out;
SharedReg959_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg959_out;
SharedReg909_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg909_out;
SharedReg809_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg809_out;
SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg954_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg472_out;
SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg660_out;
SharedReg707_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg707_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg420_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg472_out;
SharedReg956_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg956_out;
Delay8No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast <= Delay8No38_out;
SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg336_out;
SharedReg743_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg743_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg473_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg539_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg23_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg708_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg712_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg742_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg959_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg909_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg809_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg474_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg707_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg472_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg956_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay8No38_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg336_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg743_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg422_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg660_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1108_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1107_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No150_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg347_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg347_out;
SharedReg713_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg713_out;
SharedReg911_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg911_out;
SharedReg558_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg558_out;
SharedReg955_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg955_out;
SharedReg910_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg910_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg426_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg426_out;
SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg909_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg7_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg426_out;
Delay6No93_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast <= Delay6No93_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg426_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg478_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg478_out;
SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg747_out;
SharedReg823_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg823_out;
SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg747_out;
SharedReg428_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg428_out;
SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg425_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg478_out;
SharedReg481_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg481_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg478_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay6No93_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg713_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg823_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg747_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg428_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg425_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg481_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg478_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg911_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg558_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg955_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg910_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg426_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg909_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No150_out);

Delay8No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= Delay8No39_out;
SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg348_out;
SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg714_out;
SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg426_out;
SharedReg553_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg553_out;
SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg427_out;
SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg427_out;
SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg665_out;
SharedReg911_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg911_out;
SharedReg910_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg910_out;
SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg23_out;
SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg714_out;
SharedReg718_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg718_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg478_out;
SharedReg747_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg747_out;
SharedReg919_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg919_out;
SharedReg900_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg900_out;
SharedReg822_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg822_out;
SharedReg914_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg914_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg478_out;
SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg665_out;
SharedReg713_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg713_out;
SharedReg425_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg425_out;
SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg478_out;
SharedReg916_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg916_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No39_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg23_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg718_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg747_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg919_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg900_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg714_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg822_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg914_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg713_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg425_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg478_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg916_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg426_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg553_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg427_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg665_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg911_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg910_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No152_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg430_out;
SharedReg487_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg487_out;
SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg430_out;
SharedReg913_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg359_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg359_out;
SharedReg719_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg719_out;
SharedReg902_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg902_out;
SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg572_out;
SharedReg915_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg915_out;
SharedReg901_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg901_out;
SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg431_out;
SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg431_out;
SharedReg900_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg900_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg7_out;
SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg431_out;
Delay6No94_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast <= Delay6No94_out;
SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg431_out;
SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg484_out;
SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg484_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg753_out;
SharedReg836_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg836_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg753_out;
SharedReg433_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg433_out;
SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg430_out;
SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg430_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg487_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg900_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay6No94_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg431_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg484_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg836_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg753_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg433_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg430_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg913_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg359_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg719_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg902_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg572_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg915_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg901_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No152_out);

SharedReg900_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg430_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg430_out;
SharedReg906_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg725_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg725_out;
SharedReg360_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg360_out;
SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg720_out;
SharedReg431_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg431_out;
SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg432_out;
SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg432_out;
SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg670_out;
SharedReg902_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg902_out;
SharedReg901_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg901_out;
SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg23_out;
SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg720_out;
SharedReg724_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg724_out;
SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg484_out;
SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg753_out;
Delay9No31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast <= Delay9No31_out;
SharedReg453_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg453_out;
SharedReg835_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg835_out;
SharedReg904_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg904_out;
SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg484_out;
SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg670_out;
SharedReg719_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg719_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg430_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg902_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg901_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg23_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg724_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg906_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg753_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay9No31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg453_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg835_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg904_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg484_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg670_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg719_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg725_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg360_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg431_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg432_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Subtract2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_5_impl_out,
                 X => Delay1No154_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg438_out;
SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg453_out;
SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg453_out;
SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg453_out;
SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg438_out;
SharedReg435_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg435_out;
SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg903_out;
SharedReg371_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg371_out;
SharedReg759_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg759_out;
SharedReg455_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg455_out;
SharedReg586_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg586_out;
SharedReg905_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg905_out;
SharedReg454_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg454_out;
SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg436_out;
SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg436_out;
SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg453_out;
SharedReg_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg7_out;
SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg436_out;
Delay6No95_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast <= Delay6No95_out;
SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg436_out;
SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg490_out;
SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg490_out;
SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg932_out;
SharedReg849_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg849_out;
SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg932_out;
   MUX_Subtract2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg586_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg905_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg454_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg7_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay6No95_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg436_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg490_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg849_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg932_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg453_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg438_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg435_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg371_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg759_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg455_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_5_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_0_out,
                 Y => Delay1No154_out);

SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg435_out;
SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg675_out;
SharedReg673_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg673_out;
SharedReg903_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg435_out;
SharedReg935_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg935_out;
SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg765_out;
SharedReg372_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg372_out;
SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg760_out;
SharedReg436_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg436_out;
SharedReg581_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg581_out;
SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg437_out;
SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg437_out;
SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg675_out;
SharedReg455_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg455_out;
SharedReg454_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg454_out;
SharedReg16_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg23_out;
SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg760_out;
SharedReg764_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg764_out;
SharedReg490_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg490_out;
SharedReg932_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg932_out;
Delay9No32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast <= Delay9No32_out;
SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg440_out;
SharedReg848_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg848_out;
SharedReg457_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg457_out;
   MUX_Subtract2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg581_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg437_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg675_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg455_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg454_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg16_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg20_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg23_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg673_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg764_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg490_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg932_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay9No32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg848_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg457_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg903_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg435_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg765_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg372_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg760_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg436_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_5_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Subtract2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_6_impl_out,
                 X => Delay1No156_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg862_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg443_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg443_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg440_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg440_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg440_out;
SharedReg499_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg499_out;
SharedReg496_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg496_out;
SharedReg456_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg456_out;
SharedReg383_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg383_out;
SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg920_out;
SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg442_out;
SharedReg600_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg600_out;
SharedReg458_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg458_out;
SharedReg441_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg441_out;
SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg497_out;
SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg497_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg440_out;
SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg7_out;
SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg497_out;
SharedReg501_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg501_out;
SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg497_out;
SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg678_out;
SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg678_out;
   MUX_Subtract2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg383_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg600_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg458_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg441_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg920_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg4_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg7_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg501_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg497_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg678_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg443_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg440_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg499_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg496_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg456_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_6_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_0_out,
                 Y => Delay1No156_out);

SharedReg444_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg444_out;
SharedReg861_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg861_out;
SharedReg961_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg961_out;
SharedReg440_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg440_out;
SharedReg680_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg680_out;
SharedReg766_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg766_out;
SharedReg456_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg456_out;
SharedReg496_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg496_out;
SharedReg963_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg963_out;
Delay8No42_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast <= Delay8No42_out;
SharedReg384_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg384_out;
SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg921_out;
SharedReg497_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg497_out;
SharedReg595_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg595_out;
SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg498_out;
SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg498_out;
SharedReg768_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg768_out;
SharedReg442_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg442_out;
SharedReg441_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg441_out;
SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg23_out;
SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg921_out;
SharedReg925_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg925_out;
SharedReg678_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg678_out;
SharedReg960_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg960_out;
Delay9No33_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast <= Delay9No33_out;
   MUX_Subtract2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg444_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg861_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg384_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg497_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg595_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg498_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg768_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg442_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg441_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg961_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg22_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg23_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg921_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg925_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg678_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg960_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay9No33_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg440_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg680_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg766_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg456_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg496_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg963_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay8No42_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_6_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Subtract2_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_7_impl_out,
                 X => Delay1No158_out_to_Subtract2_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Subtract2_7_impl_parent_implementedSystem_port_1_cast);

SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg643_out;
SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg642_out;
SharedReg772_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg772_out;
SharedReg875_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg875_out;
SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg926_out;
SharedReg447_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg447_out;
SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg502_out;
SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg502_out;
SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg502_out;
SharedReg645_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg645_out;
SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg642_out;
SharedReg444_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg444_out;
SharedReg395_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg395_out;
SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg926_out;
SharedReg504_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg504_out;
SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg614_out;
SharedReg446_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg446_out;
SharedReg503_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg503_out;
SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg643_out;
SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg643_out;
SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg502_out;
SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg4_out;
SharedReg6_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg7_out;
SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg643_out;
SharedReg647_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg647_out;
   MUX_Subtract2_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg645_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg444_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg395_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg504_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg614_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg446_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg503_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg642_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg4_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg6_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg7_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg643_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg647_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg772_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg875_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg926_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg447_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg502_out_to_MUX_Subtract2_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_7_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_7_impl_0_out,
                 Y => Delay1No158_out);

SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg642_out;
SharedReg926_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg926_out;
Delay9No34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast <= Delay9No34_out;
SharedReg966_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg966_out;
SharedReg874_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg874_out;
SharedReg967_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg967_out;
SharedReg502_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg502_out;
SharedReg685_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg685_out;
SharedReg772_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg772_out;
SharedReg444_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg444_out;
SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg642_out;
SharedReg969_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg969_out;
Delay8No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast <= Delay8No43_out;
SharedReg396_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg396_out;
SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg927_out;
SharedReg643_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg643_out;
SharedReg609_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg609_out;
SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg644_out;
SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg644_out;
SharedReg774_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg774_out;
SharedReg504_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg504_out;
SharedReg503_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg503_out;
SharedReg16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg20_out;
SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg23_out;
SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg927_out;
SharedReg931_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg931_out;
   MUX_Subtract2_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg642_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg969_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay8No43_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg396_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg643_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg609_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg644_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg774_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay9No34_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg504_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg503_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg16_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg20_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg22_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg23_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg927_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg931_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg966_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg874_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg967_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg502_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg685_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg772_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg444_out_to_MUX_Subtract2_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_7_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_7_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Subtract2_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_8_impl_out,
                 X => Delay1No160_out_to_Subtract2_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Subtract2_8_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg451_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg510_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg510_out;
SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg638_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg505_out;
SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg450_out;
SharedReg778_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg778_out;
SharedReg888_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg888_out;
SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg726_out;
Delay4No233_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast <= Delay4No233_out;
SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg450_out;
SharedReg637_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg637_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg505_out;
SharedReg508_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg508_out;
SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg450_out;
SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg450_out;
SharedReg407_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg407_out;
SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg726_out;
SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg452_out;
SharedReg628_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg628_out;
SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg452_out;
SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg638_out;
SharedReg690_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg690_out;
SharedReg506_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg506_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg505_out;
SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg_out;
SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg4_out;
   MUX_Subtract2_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No233_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg637_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg508_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg407_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg451_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg628_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg452_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg690_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg506_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg4_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg510_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg638_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg505_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg450_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg778_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg888_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg726_out_to_MUX_Subtract2_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_8_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_8_impl_0_out,
                 Y => Delay1No160_out);

SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg23_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg727_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg727_out;
Delay6No125_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast <= Delay6No125_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg505_out;
SharedReg778_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg778_out;
SharedReg984_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg984_out;
SharedReg979_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg979_out;
SharedReg887_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg887_out;
SharedReg973_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg973_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg505_out;
SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg507_out;
SharedReg689_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg689_out;
SharedReg450_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg450_out;
SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg505_out;
SharedReg781_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg781_out;
Delay8No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast <= Delay8No44_out;
SharedReg408_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg408_out;
SharedReg779_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg779_out;
SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg451_out;
SharedReg623_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg623_out;
SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg691_out;
SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg507_out;
SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg691_out;
SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg507_out;
SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg451_out;
SharedReg16_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg16_out;
SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg20_out;
   MUX_Subtract2_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg689_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg450_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg781_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay8No44_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg408_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg779_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg727_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg623_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg691_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg507_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg451_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg16_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg20_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay6No125_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg505_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg778_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg984_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg979_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg973_out_to_MUX_Subtract2_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract2_8_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_8_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product12_8_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product12_8_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product12_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_8_impl_out,
                 X => Delay1No162_out_to_Product12_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product12_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1183_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1288_out;
SharedReg1226_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1226_out;
SharedReg389_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
SharedReg1187_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1187_out;
SharedReg1184_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1184_out;
SharedReg1189_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1218_out;
SharedReg1249_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1249_out;
SharedReg1166_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1166_out;
SharedReg1263_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1263_out;
SharedReg1278_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1278_out;
SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg876_out;
SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1168_out;
SharedReg1201_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1201_out;
SharedReg1169_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1169_out;
SharedReg1173_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1173_out;
SharedReg1204_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1204_out;
SharedReg1076_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1076_out;
SharedReg1279_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1245_out;
SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg876_out;
SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg876_out;
SharedReg1281_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1259_out;
SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1168_out;
SharedReg1196_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1196_out;
   MUX_Product12_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1183_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1288_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1263_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1278_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1201_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1169_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1173_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1204_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1076_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1279_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1226_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1244_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1245_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg876_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1281_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1259_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1168_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1196_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1187_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1184_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1189_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1218_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1249_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1166_out_to_MUX_Product12_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_8_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_8_impl_0_out,
                 Y => Delay1No162_out);

SharedReg276_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg276_out;
SharedReg1078_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1078_out;
SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg1214_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1214_out;
SharedReg614_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg614_out;
SharedReg400_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg391_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg391_out;
SharedReg86_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg86_out;
SharedReg889_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg889_out;
SharedReg1262_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1262_out;
SharedReg1077_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1077_out;
SharedReg1094_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1094_out;
SharedReg1265_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1231_out;
SharedReg290_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg290_out;
SharedReg1233_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1237_out;
SharedReg89_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg89_out;
SharedReg1219_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1219_out;
SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1076_out;
SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1076_out;
SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1076_out;
SharedReg1280_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1223_out;
SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1168_out;
SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1168_out;
SharedReg1260_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1260_out;
SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg90_out;
   MUX_Product12_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg276_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1078_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1077_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1094_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1265_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1231_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg290_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1233_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1237_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg89_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1219_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1076_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1280_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1223_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1168_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1260_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg90_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1214_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg614_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg391_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg86_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg889_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1262_out_to_MUX_Product12_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product12_8_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_8_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product22_7_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product22_7_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product22_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_7_impl_out,
                 X => Delay1No164_out_to_Product22_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product22_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1271_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1271_out;
SharedReg1212_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1212_out;
SharedReg1239_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1239_out;
SharedReg1267_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1267_out;
SharedReg1249_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1249_out;
SharedReg1247_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1247_out;
SharedReg1171_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1171_out;
SharedReg1190_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1252_out;
SharedReg1227_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1227_out;
SharedReg277_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg277_out;
SharedReg81_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg81_out;
SharedReg165_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg165_out;
SharedReg1231_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1231_out;
SharedReg1205_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1194_out;
SharedReg1242_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1196_out;
SharedReg168_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg168_out;
SharedReg1198_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1210_out;
   MUX_Product22_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1271_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1212_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg277_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg81_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg165_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1231_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1205_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1206_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1209_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1235_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1191_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1192_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1239_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1193_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1194_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1242_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1196_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg168_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1198_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1199_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1210_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1267_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1249_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1247_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1171_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1190_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1252_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1227_out_to_MUX_Product22_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product22_7_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_7_impl_0_out,
                 Y => Delay1No164_out);

SharedReg1076_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1076_out;
SharedReg278_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg278_out;
SharedReg611_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg611_out;
SharedReg1078_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1078_out;
SharedReg877_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg877_out;
SharedReg612_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg612_out;
SharedReg1270_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1270_out;
SharedReg280_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg280_out;
SharedReg1086_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
SharedReg165_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg165_out;
SharedReg1228_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1228_out;
SharedReg1229_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1229_out;
SharedReg1230_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1230_out;
SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg82_out;
SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg82_out;
SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg167_out;
SharedReg173_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg173_out;
SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg81_out;
SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg81_out;
SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg81_out;
SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg276_out;
SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg276_out;
SharedReg1168_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1168_out;
SharedReg83_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg83_out;
SharedReg1224_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1224_out;
SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg167_out;
SharedReg882_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg882_out;
SharedReg609_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg609_out;
   MUX_Product22_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1076_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg278_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1228_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1229_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1230_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg82_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg173_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg81_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg611_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg276_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1168_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg83_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1224_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg167_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg882_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg609_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1078_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg877_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg612_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1270_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg280_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg165_out_to_MUX_Product22_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product22_7_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_7_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No166_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1222_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1282_out;
SharedReg304_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg304_out;
SharedReg1239_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1258_out;
SharedReg1247_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1218_out;
SharedReg1252_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1254_out;
SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg32_out;
SharedReg1203_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1204_out;
SharedReg1205_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1233_out;
SharedReg103_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg103_out;
SharedReg1207_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1221_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1222_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1195_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1269_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1258_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1247_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1189_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1218_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1252_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1200_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1254_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1203_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1196_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1204_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1205_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1233_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg103_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1207_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1219_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1221_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1197_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1198_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1226_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1210_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1282_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg304_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1239_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No166_out);

SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg97_out;
SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg513_out;
SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg34_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg791_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg791_out;
SharedReg511_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg511_out;
SharedReg1110_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1110_out;
SharedReg1212_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1212_out;
SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg987_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg987_out;
SharedReg785_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg785_out;
SharedReg514_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg514_out;
SharedReg99_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg99_out;
SharedReg189_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg189_out;
SharedReg995_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg995_out;
SharedReg302_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg302_out;
SharedReg512_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg512_out;
SharedReg1229_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1229_out;
SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg33_out;
SharedReg186_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg186_out;
SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg33_out;
SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg97_out;
SharedReg1237_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1237_out;
SharedReg1111_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1111_out;
SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg32_out;
SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg185_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg987_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg514_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg99_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg189_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg995_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg302_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg512_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1229_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg186_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg33_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg97_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1237_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1111_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg185_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg791_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg511_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1110_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1212_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No168_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1219_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1282_out;
SharedReg316_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg316_out;
SharedReg1239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1258_out;
SharedReg1247_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1218_out;
SharedReg1252_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1254_out;
SharedReg39_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg39_out;
SharedReg1203_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1232_out;
SharedReg1206_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1207_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1219_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1220_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1282_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg316_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1269_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1258_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1247_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1189_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1218_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1252_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1200_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1221_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1254_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg39_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1203_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1204_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1232_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1206_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1209_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1207_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1222_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1195_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1196_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1197_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1198_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1226_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1210_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No168_out);

SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg107_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg107_out;
SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg527_out;
SharedReg43_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg43_out;
SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg804_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg804_out;
SharedReg525_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg525_out;
SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1118_out;
SharedReg1212_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1212_out;
SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg527_out;
SharedReg1000_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1000_out;
SharedReg798_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg798_out;
SharedReg528_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg528_out;
SharedReg109_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg109_out;
SharedReg202_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg202_out;
SharedReg1008_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1008_out;
SharedReg314_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg314_out;
SharedReg526_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg526_out;
SharedReg1229_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1229_out;
SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg40_out;
SharedReg199_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg199_out;
SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg40_out;
SharedReg1120_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1120_out;
SharedReg1010_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1010_out;
SharedReg1002_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1002_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1212_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1000_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg798_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg528_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg109_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg202_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1008_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg314_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg526_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1229_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg199_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1120_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1010_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1002_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg198_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg107_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg43_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg804_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg525_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No170_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1206_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1282_out;
SharedReg328_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg328_out;
SharedReg1239_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1258_out;
SharedReg1247_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1218_out;
SharedReg1252_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1256_out;
SharedReg212_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg212_out;
SharedReg1205_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1205_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1206_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1209_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1198_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1226_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1210_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1282_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg328_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1239_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1258_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1247_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1189_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1207_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1218_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1252_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1200_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1254_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1255_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1256_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg212_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1205_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1219_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1220_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1221_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1222_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1195_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1196_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1197_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No170_out);

SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1128_out;
SharedReg1023_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1023_out;
SharedReg1015_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1015_out;
SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg46_out;
SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg46_out;
SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg211_out;
SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg211_out;
SharedReg117_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg117_out;
SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg541_out;
SharedReg50_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg50_out;
SharedReg48_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg817_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg817_out;
SharedReg539_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg539_out;
SharedReg1126_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1126_out;
SharedReg1212_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1212_out;
SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg541_out;
SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1013_out;
SharedReg811_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg811_out;
SharedReg542_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg542_out;
SharedReg119_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg119_out;
SharedReg215_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg215_out;
SharedReg1021_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1021_out;
SharedReg326_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg326_out;
SharedReg540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg540_out;
SharedReg1012_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1012_out;
SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1128_out;
SharedReg1231_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1231_out;
SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1013_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1023_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg817_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg539_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1126_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1212_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg811_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg542_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg119_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1015_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg215_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1021_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg326_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg540_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1012_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1128_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1231_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg46_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg211_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg117_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg541_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg50_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No172_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1256_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1256_out;
SharedReg225_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg225_out;
SharedReg1205_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1282_out;
SharedReg340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg340_out;
SharedReg1239_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1258_out;
SharedReg1247_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1264_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1256_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg225_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1195_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1196_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1197_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1198_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1226_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1210_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1282_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg340_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1239_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1269_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1205_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1258_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1247_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1189_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1218_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1261_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1227_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1263_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1264_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1206_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1209_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1207_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1219_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1220_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1222_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No172_out);

SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1231_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1231_out;
SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1026_out;
SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1136_out;
SharedReg1036_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1036_out;
SharedReg1028_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg53_out;
SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg53_out;
SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg224_out;
SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg224_out;
SharedReg127_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg555_out;
SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg57_out;
SharedReg55_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg55_out;
SharedReg830_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg830_out;
SharedReg553_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg553_out;
SharedReg1134_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1134_out;
SharedReg1212_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1212_out;
SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg555_out;
SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1026_out;
SharedReg824_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg824_out;
SharedReg556_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg556_out;
SharedReg129_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg129_out;
SharedReg228_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg228_out;
SharedReg1033_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1033_out;
SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg53_out;
SharedReg554_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg554_out;
SharedReg1025_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1025_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1231_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg57_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg55_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg830_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg553_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1134_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1212_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg555_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1026_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg824_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg556_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg129_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg228_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1033_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg554_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1025_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1136_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1036_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg53_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg224_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No174_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1227_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg1256_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1256_out;
SharedReg238_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg238_out;
SharedReg1205_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1282_out;
SharedReg352_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg352_out;
SharedReg1239_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1258_out;
SharedReg1248_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1248_out;
SharedReg139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg139_out;
SharedReg1190_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1190_out;
SharedReg1047_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1047_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1227_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1220_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1221_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1222_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1195_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1196_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1197_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1198_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1226_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1210_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1282_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg352_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1239_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1269_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1258_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1248_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1190_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1047_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1256_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg238_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1205_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1206_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1209_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1207_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1219_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No174_out);

SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg568_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg1038_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1038_out;
SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1144_out;
SharedReg1231_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1231_out;
SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1039_out;
SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1144_out;
SharedReg1049_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1049_out;
SharedReg1041_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1041_out;
SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg60_out;
SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg60_out;
SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg237_out;
SharedReg137_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg137_out;
SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg569_out;
SharedReg64_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg64_out;
SharedReg62_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg62_out;
SharedReg843_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg843_out;
SharedReg567_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg567_out;
SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1142_out;
SharedReg1212_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1212_out;
SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg569_out;
SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1039_out;
SharedReg837_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg837_out;
SharedReg571_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg571_out;
SharedReg1217_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1217_out;
SharedReg242_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg242_out;
SharedReg1261_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1261_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg237_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg137_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg64_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg62_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg843_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg567_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1038_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1212_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg569_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg837_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg571_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1217_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg242_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1261_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1231_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1039_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1144_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1049_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1041_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg60_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product32_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_5_impl_out,
                 X => Delay1No176_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg1190_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1190_out;
SharedReg1060_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1060_out;
SharedReg1227_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1264_out;
SharedReg1256_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg251_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg251_out;
SharedReg1205_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1226_out;
SharedReg1210_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1282_out;
SharedReg364_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg364_out;
SharedReg1243_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1283_out;
SharedReg851_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg851_out;
SharedReg1188_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1188_out;
   MUX_Product32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1190_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1209_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1207_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1219_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1220_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1221_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1222_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1195_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1196_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1197_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1060_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1226_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1210_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1282_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg364_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1243_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1283_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg851_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1188_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1227_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1263_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1264_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg251_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1205_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1206_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_5_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_0_out,
                 Y => Delay1No176_out);

SharedReg1217_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1217_out;
SharedReg255_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg255_out;
SharedReg1261_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1261_out;
SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg67_out;
SharedReg582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg582_out;
SharedReg1051_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1051_out;
SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1152_out;
SharedReg1231_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1231_out;
SharedReg1052_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1052_out;
SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1152_out;
SharedReg1062_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1062_out;
SharedReg1054_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1054_out;
SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg67_out;
SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg67_out;
SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg250_out;
SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg250_out;
SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg147_out;
SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg583_out;
SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg71_out;
SharedReg69_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg69_out;
SharedReg856_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg856_out;
SharedReg581_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg581_out;
SharedReg1150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1150_out;
SharedReg1212_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1212_out;
SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg583_out;
SharedReg1151_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1151_out;
SharedReg1258_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1258_out;
SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg71_out;
   MUX_Product32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1217_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1062_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1054_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg250_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg69_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1261_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg856_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg581_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1212_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg583_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1151_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1258_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg71_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg67_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg582_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1051_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1231_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1052_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1152_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_5_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product32_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_6_impl_out,
                 X => Delay1No178_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1269_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1258_out;
SharedReg1248_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1248_out;
SharedReg1189_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1261_out;
SharedReg1200_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1255_out;
SharedReg1203_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1233_out;
SharedReg163_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg163_out;
SharedReg1207_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1194_out;
SharedReg1160_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1160_out;
SharedReg1223_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1223_out;
SharedReg158_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg158_out;
SharedReg1198_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1282_out;
SharedReg376_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg376_out;
SharedReg1243_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1243_out;
   MUX_Product32_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1269_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1258_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1204_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1232_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1233_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg163_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1207_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1192_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1160_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1248_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1223_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg158_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1198_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1199_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1210_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1282_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg376_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1243_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1189_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1218_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1261_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1200_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1254_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1255_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1203_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_6_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_0_out,
                 Y => Delay1No178_out);

SharedReg1065_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1065_out;
SharedReg863_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg863_out;
SharedReg599_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg599_out;
SharedReg159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg267_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg267_out;
SharedReg1072_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1072_out;
SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg374_out;
SharedReg596_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg596_out;
SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1064_out;
SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg75_out;
SharedReg264_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg264_out;
SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg75_out;
SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg157_out;
SharedReg1237_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1237_out;
SharedReg1159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1159_out;
SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg155_out;
SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg155_out;
SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg374_out;
SharedReg1246_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1246_out;
SharedReg76_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg76_out;
SharedReg1224_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1224_out;
SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg157_out;
SharedReg869_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg869_out;
SharedReg595_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg595_out;
SharedReg1158_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1158_out;
SharedReg1212_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1212_out;
SharedReg597_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg597_out;
   MUX_Product32_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1065_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg863_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg264_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1237_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg155_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1246_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg599_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg76_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1224_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg157_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg869_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg595_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1158_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1212_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg597_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1072_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg374_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg596_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg75_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_6_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product32_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_7_impl_out,
                 X => Delay1No180_out_to_Product32_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product32_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1282_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1282_out;
SharedReg388_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg1243_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1243_out;
SharedReg1269_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1269_out;
SharedReg1258_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1258_out;
SharedReg1248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1248_out;
SharedReg1189_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1261_out;
SharedReg1200_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1200_out;
SharedReg1254_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1255_out;
SharedReg1203_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1204_out;
SharedReg1232_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1233_out;
SharedReg173_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg173_out;
SharedReg1207_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1207_out;
SharedReg1191_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1192_out;
SharedReg1193_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1193_out;
SharedReg1194_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1194_out;
SharedReg1168_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1168_out;
SharedReg1223_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1223_out;
SharedReg1197_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1226_out;
SharedReg874_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg874_out;
   MUX_Product32_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1282_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1254_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1255_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1203_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1204_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1232_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1233_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg173_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1207_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1191_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1192_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1243_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1193_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1194_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1168_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1223_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1197_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1198_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1226_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg874_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1269_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1258_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1248_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1189_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1218_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1261_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1200_out_to_MUX_Product32_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_7_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_7_impl_0_out,
                 Y => Delay1No180_out);

SharedReg1166_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1166_out;
SharedReg1212_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1212_out;
SharedReg611_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg611_out;
SharedReg1078_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1078_out;
SharedReg876_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg876_out;
SharedReg613_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg613_out;
SharedReg169_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg169_out;
SharedReg280_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg280_out;
SharedReg1085_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1085_out;
SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg386_out;
SharedReg610_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg610_out;
SharedReg1077_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1077_out;
SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg82_out;
SharedReg277_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg277_out;
SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg82_out;
SharedReg167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg167_out;
SharedReg1237_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1237_out;
SharedReg1167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1167_out;
SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg165_out;
SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg165_out;
SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg386_out;
SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg386_out;
SharedReg1246_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1246_out;
SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg83_out;
SharedReg85_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg85_out;
SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg83_out;
SharedReg882_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg882_out;
SharedReg1210_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1210_out;
   MUX_Product32_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1166_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1212_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg610_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1077_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg277_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg82_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1237_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1167_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg165_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg611_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1246_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg85_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg83_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg882_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1210_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1078_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg876_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg613_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg169_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg280_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1085_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg386_out_to_MUX_Product32_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product32_7_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_7_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product6_8_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product6_8_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product6_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_8_impl_out,
                 X => Delay1No182_out_to_Product6_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product6_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1197_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1198_out;
SharedReg1199_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1199_out;
SharedReg1210_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1210_out;
SharedReg1282_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1282_out;
SharedReg1090_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1090_out;
SharedReg1239_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1239_out;
SharedReg1269_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1269_out;
SharedReg890_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg890_out;
SharedReg1247_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1247_out;
SharedReg1189_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1189_out;
SharedReg1190_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1190_out;
SharedReg1252_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1252_out;
SharedReg1200_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1200_out;
SharedReg1263_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1263_out;
SharedReg88_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg88_out;
SharedReg1203_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1203_out;
SharedReg290_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg290_out;
SharedReg1205_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1233_out;
SharedReg183_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg183_out;
SharedReg1235_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1191_out;
SharedReg1192_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1192_out;
SharedReg1221_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1196_out;
   MUX_Product6_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1197_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1198_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1189_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1190_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1252_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1200_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1263_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg88_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1203_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg290_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1205_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1233_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1199_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg183_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1235_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1191_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1192_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1221_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1222_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1195_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1196_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1210_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1282_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1090_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1239_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1269_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg890_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1247_out_to_MUX_Product6_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_8_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_8_impl_0_out,
                 Y => Delay1No182_out);

SharedReg92_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg90_out;
SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg623_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg623_out;
SharedReg1174_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1174_out;
SharedReg1277_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1277_out;
SharedReg625_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg625_out;
SharedReg1091_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1091_out;
SharedReg1258_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1258_out;
SharedReg626_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg626_out;
SharedReg179_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg179_out;
SharedReg294_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg294_out;
SharedReg1099_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1099_out;
SharedReg398_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg398_out;
SharedReg624_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg624_out;
SharedReg1229_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1229_out;
SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg89_out;
SharedReg1231_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1231_out;
SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg89_out;
SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg177_out;
SharedReg1237_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1237_out;
SharedReg88_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg88_out;
SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg175_out;
SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg175_out;
SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg289_out;
SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg289_out;
SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg177_out;
SharedReg889_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg889_out;
   MUX_Product6_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg179_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg294_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1099_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg398_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg624_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1229_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1231_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg89_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1237_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg88_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg175_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg289_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg177_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg889_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg623_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1174_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1277_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg625_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1091_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1258_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg626_out_to_MUX_Product6_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product6_8_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_8_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product23_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_0_impl_out,
                 X => Delay1No184_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg1242_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1199_out;
SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg783_out;
SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1110_out;
SharedReg986_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg986_out;
SharedReg1243_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1283_out;
SharedReg786_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg786_out;
SharedReg1248_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1248_out;
SharedReg99_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg99_out;
SharedReg1190_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1190_out;
SharedReg1261_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1263_out;
SharedReg1255_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1256_out;
SharedReg186_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg186_out;
SharedReg1232_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1232_out;
SharedReg1206_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1207_out;
SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg95_out;
SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg302_out;
   MUX_Product23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1242_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1283_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg786_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1248_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg99_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1190_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1261_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1227_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1263_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1255_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1256_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1196_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg186_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1232_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1206_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1209_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1207_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg302_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1224_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1225_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1199_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg986_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1243_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_0_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_0_out,
                 Y => Delay1No184_out);

SharedReg1222_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1222_out;
SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1111_out;
SharedReg785_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg785_out;
SharedReg36_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg34_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg34_out;
SharedReg1210_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1277_out;
SharedReg513_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1111_out;
SharedReg1258_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1258_out;
SharedReg515_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg515_out;
SharedReg1217_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1217_out;
SharedReg190_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg190_out;
SharedReg994_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg994_out;
SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg32_out;
SharedReg512_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg512_out;
SharedReg986_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg986_out;
SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1112_out;
SharedReg1231_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1231_out;
SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg33_out;
SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1112_out;
SharedReg997_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg997_out;
SharedReg989_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg989_out;
SharedReg1219_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1221_out;
   MUX_Product23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1222_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1111_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1258_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg515_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1217_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg190_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg994_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg512_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg986_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg785_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1231_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg33_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1112_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg997_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg989_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1219_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1220_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1221_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg34_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1210_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1284_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1277_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_0_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product23_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_1_impl_out,
                 X => Delay1No186_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg314_out;
SharedReg1242_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1199_out;
SharedReg796_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg796_out;
SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1118_out;
SharedReg999_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg999_out;
SharedReg1243_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1283_out;
SharedReg799_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg799_out;
SharedReg1248_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1248_out;
SharedReg109_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg109_out;
SharedReg1190_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1190_out;
SharedReg1261_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1263_out;
SharedReg1255_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1256_out;
SharedReg199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg199_out;
SharedReg1205_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1235_out;
   MUX_Product23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg999_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1243_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1283_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg799_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1248_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg109_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1190_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1261_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1227_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1263_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1255_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1256_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1205_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1206_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1209_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1235_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg314_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1242_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1196_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1224_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1225_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1199_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg796_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_1_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_0_out,
                 Y => Delay1No186_out);

SharedReg1219_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1222_out;
SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1119_out;
SharedReg798_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg798_out;
SharedReg43_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg43_out;
SharedReg107_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg107_out;
SharedReg41_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg41_out;
SharedReg1210_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1277_out;
SharedReg527_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg527_out;
SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1119_out;
SharedReg1258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1258_out;
SharedReg529_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg529_out;
SharedReg1217_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1217_out;
SharedReg203_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg203_out;
SharedReg1007_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1007_out;
SharedReg39_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg39_out;
SharedReg526_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg526_out;
SharedReg999_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg999_out;
SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1120_out;
SharedReg1231_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1231_out;
SharedReg1000_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1000_out;
SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1121_out;
SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1125_out;
SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1119_out;
   MUX_Product23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1219_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1220_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1284_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1277_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg527_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1258_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg529_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1217_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg203_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1007_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg39_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1221_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg526_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg999_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1231_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1000_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1222_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg798_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg43_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg107_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg41_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1210_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_1_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product23_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_2_impl_out,
                 X => Delay1No188_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1206_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1235_out;
SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg115_out;
SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg326_out;
SharedReg1242_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1199_out;
SharedReg809_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg809_out;
SharedReg1126_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1126_out;
SharedReg1012_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1012_out;
SharedReg1243_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1283_out;
SharedReg812_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg812_out;
SharedReg1248_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1248_out;
SharedReg119_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg119_out;
SharedReg1190_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1190_out;
SharedReg1261_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1264_out;
SharedReg1128_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1128_out;
SharedReg1257_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1205_out;
   MUX_Product23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1206_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1209_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1225_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1199_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg809_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1126_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1012_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1243_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1283_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg812_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1248_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg119_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1235_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1190_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1261_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1227_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1263_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1264_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1128_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1257_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1205_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg115_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1242_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1196_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1224_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_2_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_0_out,
                 Y => Delay1No188_out);

SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1133_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1133_out;
SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1127_out;
SharedReg1219_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1222_out;
SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1127_out;
SharedReg811_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg811_out;
SharedReg50_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg50_out;
SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg117_out;
SharedReg48_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg48_out;
SharedReg1210_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1277_out;
SharedReg541_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg541_out;
SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1127_out;
SharedReg1258_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1258_out;
SharedReg543_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg543_out;
SharedReg1217_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1217_out;
SharedReg216_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg216_out;
SharedReg1020_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1020_out;
SharedReg46_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg46_out;
SharedReg540_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg540_out;
SharedReg1012_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1012_out;
SharedReg1265_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1265_out;
SharedReg1013_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1013_out;
SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1129_out;
   MUX_Product23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1133_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg48_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1210_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1284_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1277_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg541_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1258_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg543_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1217_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg216_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1020_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg46_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg540_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1012_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1265_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1013_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1129_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1219_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1220_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1221_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1222_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1127_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg811_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg50_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_2_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product23_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_3_impl_out,
                 X => Delay1No190_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1136_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1257_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1235_out;
SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg125_out;
SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg125_out;
SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg338_out;
SharedReg1242_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1199_out;
SharedReg822_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg822_out;
SharedReg1134_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1134_out;
SharedReg1025_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1025_out;
SharedReg1243_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1283_out;
SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg825_out;
SharedReg1248_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1248_out;
SharedReg129_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg129_out;
SharedReg1190_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1190_out;
SharedReg1034_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1034_out;
SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg338_out;
SharedReg1201_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1255_out;
   MUX_Product23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1257_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1242_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1196_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1224_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1225_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1199_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg822_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1134_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1025_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1243_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1283_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1205_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1248_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg129_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1190_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1034_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1201_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1255_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1206_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1209_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1235_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg125_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg338_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_3_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_0_out,
                 Y => Delay1No190_out);

SharedReg1265_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1265_out;
SharedReg1026_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1026_out;
SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1137_out;
SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1141_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1141_out;
SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1135_out;
SharedReg1219_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1222_out;
SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1135_out;
SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg824_out;
SharedReg57_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg57_out;
SharedReg127_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
SharedReg55_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg55_out;
SharedReg1210_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1277_out;
SharedReg555_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg555_out;
SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1135_out;
SharedReg1258_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1258_out;
SharedReg557_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg557_out;
SharedReg1217_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1217_out;
SharedReg229_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg229_out;
SharedReg1261_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1227_out;
SharedReg54_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg54_out;
SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg824_out;
   MUX_Product23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1265_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1026_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg57_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg55_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1210_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1284_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1277_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg555_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1258_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg557_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1217_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg229_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1261_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1227_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg54_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg824_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1141_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1135_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1219_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1220_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1221_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1222_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_3_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product23_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_4_impl_out,
                 X => Delay1No192_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast);

SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg1201_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1255_out;
SharedReg1144_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1144_out;
SharedReg1257_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1235_out;
SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg135_out;
SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg135_out;
SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg350_out;
SharedReg1242_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1199_out;
SharedReg835_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg835_out;
SharedReg1142_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1142_out;
SharedReg1038_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1038_out;
SharedReg1243_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1283_out;
SharedReg838_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg838_out;
SharedReg1188_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1208_out;
   MUX_Product23_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1201_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg350_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1242_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1196_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1224_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1225_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1199_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg835_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1142_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1255_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1038_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1243_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1283_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg838_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1188_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1218_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1208_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1144_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1257_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1205_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1206_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1209_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1235_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg135_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_4_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_0_out,
                 Y => Delay1No192_out);

SharedReg1227_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1227_out;
SharedReg61_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg837_out;
SharedReg1265_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1265_out;
SharedReg1039_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1039_out;
SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1145_out;
SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1145_out;
SharedReg1149_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1149_out;
SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1143_out;
SharedReg1219_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1222_out;
SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1143_out;
SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg837_out;
SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg64_out;
SharedReg137_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg137_out;
SharedReg62_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg1210_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1277_out;
SharedReg569_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg569_out;
SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1143_out;
SharedReg1258_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1258_out;
SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg64_out;
SharedReg354_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg354_out;
SharedReg242_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg242_out;
SharedReg66_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg66_out;
   MUX_Product23_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1227_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1220_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1221_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1222_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg137_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1210_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1284_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg837_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1277_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg569_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1258_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg64_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg354_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg242_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg66_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1265_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1039_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1145_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1149_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1143_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1219_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_4_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product23_8_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product23_8_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product23_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_8_impl_out,
                 X => Delay1No194_out_to_Product23_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product23_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1224_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1199_out;
SharedReg887_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg887_out;
SharedReg1174_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1174_out;
SharedReg1184_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1184_out;
SharedReg1243_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1243_out;
SharedReg1283_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1283_out;
SharedReg1187_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1187_out;
SharedReg1248_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1248_out;
SharedReg179_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg179_out;
SharedReg1218_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1218_out;
SharedReg1261_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1227_out;
SharedReg1201_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1256_out;
SharedReg1257_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1257_out;
SharedReg1232_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1232_out;
SharedReg1206_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1220_out;
SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg398_out;
SharedReg1242_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1242_out;
SharedReg1223_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1223_out;
   MUX_Product23_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1224_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1225_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg179_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1218_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1261_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1227_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1201_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1255_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1256_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1257_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1232_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1206_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1199_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1209_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1207_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1219_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1220_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg398_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1242_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1223_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg887_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1174_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1184_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1243_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1283_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1187_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1248_out_to_MUX_Product23_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_8_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_8_impl_0_out,
                 Y => Delay1No194_out);

SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg177_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg177_out;
SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg1210_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1284_out;
SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg625_out;
SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1175_out;
SharedReg178_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg178_out;
SharedReg627_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg627_out;
SharedReg1217_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1217_out;
SharedReg294_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg294_out;
SharedReg1098_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1098_out;
SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg88_out;
SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg89_out;
SharedReg1090_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1090_out;
SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1176_out;
SharedReg1091_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1091_out;
SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg89_out;
SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1176_out;
SharedReg1101_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1101_out;
SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1175_out;
SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg88_out;
SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg88_out;
SharedReg1221_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1222_out;
SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1175_out;
SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg625_out;
   MUX_Product23_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg177_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1217_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg294_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1098_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1090_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1091_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1176_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg92_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1101_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg88_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1221_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1222_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1210_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1284_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg625_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1175_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg178_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg627_out_to_MUX_Product23_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product23_8_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_8_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product33_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_0_impl_out,
                 X => Delay1No196_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1241_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1223_out;
SharedReg99_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg1199_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1184_out;
SharedReg785_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg785_out;
SharedReg1285_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1218_out;
SharedReg995_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg995_out;
SharedReg302_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg302_out;
SharedReg1201_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1201_out;
SharedReg1264_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1264_out;
SharedReg1112_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1112_out;
SharedReg1257_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1240_out;
   MUX_Product33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1241_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1274_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1285_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1187_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1188_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1189_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1218_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg995_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg302_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1201_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1264_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1112_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1223_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1257_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1205_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1206_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1209_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1235_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1191_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1273_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1240_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg99_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1199_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1286_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1183_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1184_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg785_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_0_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_0_out,
                 Y => Delay1No196_out);

SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg785_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg785_out;
SharedReg513_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg513_out;
SharedReg1224_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1225_out;
SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg985_out;
SharedReg95_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg95_out;
SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg1243_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1243_out;
SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1111_out;
SharedReg98_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg98_out;
SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg36_out;
SharedReg306_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg306_out;
SharedReg190_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg190_out;
SharedReg1261_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1227_out;
SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg33_out;
SharedReg986_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg986_out;
SharedReg1265_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1265_out;
SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg987_out;
SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg987_out;
SharedReg1113_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1113_out;
SharedReg1117_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1117_out;
SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1111_out;
SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg985_out;
SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg985_out;
SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg985_out;
   MUX_Product33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg785_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg306_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg190_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1261_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1227_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg986_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1265_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg513_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg987_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1113_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1117_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1111_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1224_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1225_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg985_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg95_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1243_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_0_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product33_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_1_impl_out,
                 X => Delay1No198_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1191_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1223_out;
SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg109_out;
SharedReg41_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg1199_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1184_out;
SharedReg798_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg798_out;
SharedReg1285_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1218_out;
SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1008_out;
SharedReg314_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg314_out;
SharedReg1201_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1201_out;
SharedReg1264_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1264_out;
SharedReg1120_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1120_out;
SharedReg1257_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1237_out;
SharedReg1002_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1002_out;
   MUX_Product33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1191_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1273_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1183_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1184_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg798_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1285_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1187_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1188_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1189_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1218_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg314_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1240_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1201_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1264_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1120_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1257_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1205_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1233_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1237_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1002_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1241_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1223_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1199_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1286_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_1_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_0_out,
                 Y => Delay1No198_out);

SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg998_out;
SharedReg798_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg798_out;
SharedReg527_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg527_out;
SharedReg1224_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1225_out;
SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg43_out;
SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg998_out;
SharedReg105_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg105_out;
SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg40_out;
SharedReg1243_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1243_out;
SharedReg1119_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1119_out;
SharedReg108_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg108_out;
SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg43_out;
SharedReg318_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg318_out;
SharedReg203_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg203_out;
SharedReg1261_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1227_out;
SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg40_out;
SharedReg999_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg999_out;
SharedReg1265_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1265_out;
SharedReg1000_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1000_out;
SharedReg1121_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1121_out;
SharedReg1120_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1120_out;
SharedReg1010_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1010_out;
SharedReg1235_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1235_out;
   MUX_Product33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg105_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1243_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1119_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg108_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg318_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg203_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1261_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1227_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg40_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg999_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1265_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1000_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1121_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1120_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1010_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1235_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg798_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1224_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1225_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg43_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg998_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_1_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product33_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_2_impl_out,
                 X => Delay1No200_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1233_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1237_out;
SharedReg1015_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1015_out;
SharedReg1191_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1223_out;
SharedReg119_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg119_out;
SharedReg48_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg1199_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1184_out;
SharedReg811_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg811_out;
SharedReg1285_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1218_out;
SharedReg1021_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1021_out;
SharedReg326_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg326_out;
SharedReg1201_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1232_out;
   MUX_Product33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1233_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1237_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1199_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1286_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1183_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1184_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg811_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1285_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1187_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1188_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1189_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1015_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1218_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1021_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg326_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1201_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1255_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1256_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1266_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1232_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1191_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1273_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1240_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1241_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1274_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1223_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg119_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_2_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_0_out,
                 Y => Delay1No200_out);

SharedReg1128_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1128_out;
SharedReg1023_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1023_out;
SharedReg1235_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1235_out;
SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1011_out;
SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg811_out;
SharedReg541_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg541_out;
SharedReg1224_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1225_out;
SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg50_out;
SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1011_out;
SharedReg115_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg115_out;
SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg47_out;
SharedReg1243_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1243_out;
SharedReg1127_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1127_out;
SharedReg118_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg118_out;
SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg50_out;
SharedReg330_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg330_out;
SharedReg216_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg216_out;
SharedReg1261_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1227_out;
SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg47_out;
SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg811_out;
SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg811_out;
SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1013_out;
SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1013_out;
   MUX_Product33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1128_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1023_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1225_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg115_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1243_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1127_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg118_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg50_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg330_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1235_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg216_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1261_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1227_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg47_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1013_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1011_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg811_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg541_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1224_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_2_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product33_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_3_impl_out,
                 X => Delay1No202_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1256_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1237_out;
SharedReg1028_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg1191_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1223_out;
SharedReg129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg129_out;
SharedReg55_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg55_out;
SharedReg1199_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1184_out;
SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg824_out;
SharedReg1285_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1208_out;
SharedReg1253_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1254_out;
SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg824_out;
   MUX_Product33_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1256_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1266_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1274_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1223_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg55_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1199_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1286_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1183_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1184_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1285_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1232_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1187_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1188_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1189_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1218_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1208_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1253_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1254_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg824_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1233_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1237_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1191_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1273_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1240_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1241_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_3_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_0_out,
                 Y => Delay1No202_out);

SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg824_out;
SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1026_out;
SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1026_out;
SharedReg1136_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1136_out;
SharedReg1036_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1036_out;
SharedReg1235_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1235_out;
SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1024_out;
SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1024_out;
SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1024_out;
SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1024_out;
SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg824_out;
SharedReg555_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg555_out;
SharedReg1224_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1225_out;
SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg57_out;
SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1024_out;
SharedReg125_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg125_out;
SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg54_out;
SharedReg1243_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1243_out;
SharedReg1135_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1135_out;
SharedReg128_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg57_out;
SharedReg342_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg342_out;
SharedReg229_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg229_out;
SharedReg59_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg59_out;
SharedReg1134_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1134_out;
SharedReg1025_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1025_out;
SharedReg1264_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1264_out;
   MUX_Product33_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg824_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg555_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1224_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1225_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg125_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1243_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1135_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1026_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg57_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg342_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg229_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg59_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1134_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1025_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1264_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1136_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1036_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1235_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1024_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_3_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product33_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_4_impl_out,
                 X => Delay1No204_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1253_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1254_out;
SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg837_out;
SharedReg1256_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1237_out;
SharedReg1041_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1041_out;
SharedReg1191_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1223_out;
SharedReg139_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg139_out;
SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg62_out;
SharedReg1199_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1184_out;
SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg837_out;
SharedReg1285_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1187_out;
SharedReg1216_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1216_out;
SharedReg354_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg354_out;
SharedReg1190_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1190_out;
SharedReg1236_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1236_out;
   MUX_Product33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1253_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1254_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1273_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1240_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1241_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1274_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1223_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg139_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1199_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1286_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1183_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1184_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg837_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1285_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1187_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1216_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg354_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1190_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1236_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1256_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1266_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1232_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1233_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1237_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1041_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1191_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_4_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_0_out,
                 Y => Delay1No204_out);

SharedReg1142_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1142_out;
SharedReg1038_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1038_out;
SharedReg1264_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg837_out;
SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1039_out;
SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1039_out;
SharedReg1144_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1144_out;
SharedReg1049_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1049_out;
SharedReg1235_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1235_out;
SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1037_out;
SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1037_out;
SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1037_out;
SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1037_out;
SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg837_out;
SharedReg569_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg569_out;
SharedReg1224_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1225_out;
SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg64_out;
SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1037_out;
SharedReg135_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg135_out;
SharedReg61_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg61_out;
SharedReg1243_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1243_out;
SharedReg1143_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1143_out;
SharedReg138_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg138_out;
SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg64_out;
SharedReg1217_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1217_out;
SharedReg65_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg66_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg66_out;
   MUX_Product33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1142_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1038_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg569_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1224_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1225_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg135_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg61_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1243_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1143_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg138_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg64_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1217_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg66_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg837_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1039_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1144_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1049_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1235_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1037_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_4_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product33_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_5_impl_out,
                 X => Delay1No206_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1189_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1208_out;
SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg362_out;
SharedReg1201_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1255_out;
SharedReg1152_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1152_out;
SharedReg1257_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1235_out;
SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg145_out;
SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg145_out;
SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg362_out;
SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg362_out;
SharedReg1242_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1199_out;
SharedReg848_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg848_out;
SharedReg1150_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1150_out;
SharedReg1051_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1051_out;
SharedReg850_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg850_out;
SharedReg1285_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1187_out;
SharedReg1216_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1216_out;
   MUX_Product33_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1189_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1218_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1209_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1235_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg145_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1242_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1196_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1224_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1225_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1208_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1199_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg848_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1150_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1051_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg850_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1285_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1187_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1216_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg362_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1201_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1255_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1152_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1257_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1205_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1206_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_5_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_5_impl_0_out,
                 Y => Delay1No206_out);

SharedReg366_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg366_out;
SharedReg255_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg255_out;
SharedReg73_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg73_out;
SharedReg1227_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1227_out;
SharedReg68_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg68_out;
SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg850_out;
SharedReg1265_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1265_out;
SharedReg1052_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1052_out;
SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1153_out;
SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1153_out;
SharedReg1157_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1157_out;
SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1151_out;
SharedReg1219_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1222_out;
SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1151_out;
SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg850_out;
SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg71_out;
SharedReg147_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg147_out;
SharedReg69_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg69_out;
SharedReg1210_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1277_out;
SharedReg1243_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1243_out;
SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1151_out;
SharedReg148_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg148_out;
SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg71_out;
   MUX_Product33_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg366_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1157_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1219_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1220_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1221_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1222_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg147_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg73_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg69_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1210_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1284_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1277_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1243_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1151_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg148_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg71_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1227_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg68_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg850_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1265_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1052_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1153_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_5_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_5_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product33_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_6_impl_out,
                 X => Delay1No208_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1283_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1283_out;
SharedReg864_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg864_out;
SharedReg1188_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1188_out;
SharedReg159_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg1190_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1190_out;
SharedReg1073_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1073_out;
SharedReg1227_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg1256_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1256_out;
SharedReg264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg264_out;
SharedReg1205_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1196_out;
SharedReg1197_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1197_out;
SharedReg1198_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1198_out;
SharedReg1226_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1226_out;
SharedReg861_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg861_out;
SharedReg1158_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1158_out;
SharedReg1064_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1064_out;
SharedReg863_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg863_out;
   MUX_Product33_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1283_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg864_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1205_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1206_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1209_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1207_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1219_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1220_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1221_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1222_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1195_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1188_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1196_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1197_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1198_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1226_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg861_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1158_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1064_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg863_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1190_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1073_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1227_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1256_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_6_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_6_impl_0_out,
                 Y => Delay1No208_out);

SharedReg1159_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1159_out;
SharedReg1258_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1258_out;
SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg1217_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1217_out;
SharedReg268_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg268_out;
SharedReg1261_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1261_out;
SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg74_out;
SharedReg596_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg596_out;
SharedReg1064_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1064_out;
SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1160_out;
SharedReg1231_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1231_out;
SharedReg1065_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1065_out;
SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1160_out;
SharedReg1075_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1075_out;
SharedReg1067_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1067_out;
SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg74_out;
SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg74_out;
SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg263_out;
SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg263_out;
SharedReg157_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg157_out;
SharedReg597_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg597_out;
SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg78_out;
SharedReg76_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg76_out;
SharedReg869_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg869_out;
SharedReg1210_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1210_out;
SharedReg1284_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1277_out;
SharedReg1243_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1243_out;
   MUX_Product33_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1159_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1258_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1231_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1065_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1075_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1067_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg263_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg157_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg597_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg78_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg76_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg869_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1210_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1284_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1277_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1243_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1217_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg268_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1261_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg74_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg596_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1064_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1160_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_6_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_6_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product33_7_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product33_7_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product33_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_7_impl_out,
                 X => Delay1No210_out_to_Product33_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product33_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1166_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1166_out;
SharedReg1077_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1077_out;
SharedReg876_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg1283_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1283_out;
SharedReg877_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg877_out;
SharedReg1188_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1188_out;
SharedReg169_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg169_out;
SharedReg1190_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1190_out;
SharedReg1086_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
SharedReg1227_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1227_out;
SharedReg1263_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1264_out;
SharedReg1256_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
SharedReg277_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg277_out;
SharedReg1205_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1207_out;
SharedReg1219_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1222_out;
SharedReg1195_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1195_out;
SharedReg1196_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1286_out;
   MUX_Product33_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1166_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1077_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1263_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1264_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg277_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1205_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1206_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1209_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1207_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1219_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1220_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg876_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1221_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1222_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1195_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1196_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1224_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1225_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1199_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1286_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1283_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg877_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1188_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg169_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1190_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1227_out_to_MUX_Product33_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_7_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_7_impl_0_out,
                 Y => Delay1No210_out);

SharedReg1284_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1284_out;
SharedReg1277_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1277_out;
SharedReg1243_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1243_out;
SharedReg1167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1167_out;
SharedReg1258_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1258_out;
SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg85_out;
SharedReg1217_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1217_out;
SharedReg281_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg281_out;
SharedReg1261_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1261_out;
SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg81_out;
SharedReg610_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg610_out;
SharedReg1077_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1077_out;
SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1168_out;
SharedReg1231_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1231_out;
SharedReg1078_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1078_out;
SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1168_out;
SharedReg1088_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1088_out;
SharedReg1080_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1080_out;
SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg81_out;
SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg81_out;
SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg276_out;
SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg276_out;
SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg167_out;
SharedReg611_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg611_out;
SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg85_out;
SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg167_out;
SharedReg83_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg83_out;
SharedReg1076_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1076_out;
   MUX_Product33_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1284_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1277_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg610_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1077_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1231_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1078_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1168_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1088_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1080_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1243_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg276_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg611_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg83_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1076_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1167_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1258_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg85_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1217_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg281_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1261_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg81_out_to_MUX_Product33_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_7_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_7_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product33_8_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product33_8_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product33_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_8_impl_out,
                 X => Delay1No212_out_to_Product33_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product33_8_impl_parent_implementedSystem_port_1_cast);

SharedReg179_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg90_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg90_out;
SharedReg1251_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1183_out;
SharedReg1212_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1212_out;
SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg889_out;
SharedReg1285_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1285_out;
SharedReg178_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg178_out;
SharedReg1188_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1189_out;
SharedReg1190_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1190_out;
SharedReg1099_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1099_out;
SharedReg398_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg398_out;
SharedReg1254_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1254_out;
SharedReg1264_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1264_out;
SharedReg1176_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1176_out;
SharedReg1266_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1266_out;
SharedReg1205_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1209_out;
SharedReg1207_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1207_out;
SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg175_out;
SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg175_out;
SharedReg1240_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1274_out;
SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg889_out;
   MUX_Product33_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg90_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1189_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1190_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1099_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg398_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1254_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1264_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1176_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1266_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1205_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1206_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1251_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1209_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1207_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg175_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1240_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1241_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1274_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1286_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1183_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1212_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg889_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1285_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg178_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1188_out_to_MUX_Product33_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_8_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_8_impl_0_out,
                 Y => Delay1No212_out);

SharedReg1224_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1225_out;
SharedReg1176_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1176_out;
SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1089_out;
SharedReg175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg89_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg1243_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1243_out;
SharedReg1175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1175_out;
SharedReg1215_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1215_out;
SharedReg92_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg92_out;
SharedReg402_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg402_out;
SharedReg93_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg93_out;
SharedReg1261_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1261_out;
SharedReg1227_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1227_out;
SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1090_out;
SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1090_out;
SharedReg1265_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1265_out;
SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1091_out;
SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1091_out;
SharedReg1177_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1177_out;
SharedReg1181_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1181_out;
SharedReg1093_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1093_out;
SharedReg1219_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1220_out;
SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1089_out;
SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1089_out;
SharedReg889_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg889_out;
SharedReg1223_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1223_out;
   MUX_Product33_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1224_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1225_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg402_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg93_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1261_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1227_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1090_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1265_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1091_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1177_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1176_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1181_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1093_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1219_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1220_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg889_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1223_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1089_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg89_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1243_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1175_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1215_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg92_out_to_MUX_Product33_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product33_8_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_8_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Subtract4_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_0_impl_out,
                 X => Delay1No214_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast);

Delay10No18_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast <= Delay10No18_out;
SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg412_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg412_out;
SharedReg414_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg414_out;
SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg648_out;
SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg100_out;
SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg695_out;
SharedReg308_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg308_out;
SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg96_out;
SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg34_out;
SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg648_out;
SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg695_out;
SharedReg1102_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1102_out;
SharedReg792_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg792_out;
SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg733_out;
SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg695_out;
SharedReg460_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg460_out;
SharedReg783_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg783_out;
SharedReg939_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg939_out;
SharedReg185_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg185_out;
SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg100_out;
SharedReg697_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg697_out;
SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg733_out;
SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg733_out;
SharedReg696_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg696_out;
   MUX_Subtract4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay10No18_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg308_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg34_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1102_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg792_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg460_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg5_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg783_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg939_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg185_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg697_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg733_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg696_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg9_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg412_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg414_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg648_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg100_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg695_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_0_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_0_out,
                 Y => Delay1No214_out);

SharedReg649_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg649_out;
SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg697_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg697_out;
SharedReg699_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg699_out;
SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg732_out;
SharedReg193_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg193_out;
SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg411_out;
SharedReg310_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg310_out;
SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg185_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg185_out;
SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg732_out;
SharedReg698_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg698_out;
SharedReg700_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg700_out;
SharedReg524_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg524_out;
SharedReg695_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg695_out;
SharedReg940_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg940_out;
SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg732_out;
SharedReg511_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg511_out;
SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1103_out;
SharedReg302_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg302_out;
SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg95_out;
SharedReg733_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg733_out;
SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1104_out;
SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1104_out;
SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1103_out;
   MUX_Subtract4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg649_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg310_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg185_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg698_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg700_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg524_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg695_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg940_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg511_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg302_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg95_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg733_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1104_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1103_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg25_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg697_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg699_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg732_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg193_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_0_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No216_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg738_out;
SharedReg702_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg702_out;
SharedReg654_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg654_out;
Delay10No19_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= Delay10No19_out;
SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg417_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg417_out;
SharedReg419_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg419_out;
SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg653_out;
SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg110_out;
SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg701_out;
SharedReg320_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg320_out;
SharedReg106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg106_out;
SharedReg41_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg41_out;
SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg653_out;
SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg701_out;
SharedReg1106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1106_out;
SharedReg805_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg805_out;
SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg738_out;
SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg701_out;
SharedReg466_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg466_out;
SharedReg796_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg796_out;
SharedReg946_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg946_out;
SharedReg198_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg198_out;
SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg110_out;
SharedReg703_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg703_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg702_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg320_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg41_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg653_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1106_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg805_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg654_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg738_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg701_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg466_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg796_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg946_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg198_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg110_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg703_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay10No19_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg9_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg417_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg419_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No216_out);

SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1108_out;
SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg947_out;
SharedReg467_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg467_out;
SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg703_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg703_out;
SharedReg705_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg705_out;
SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg737_out;
SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg206_out;
SharedReg416_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg416_out;
SharedReg322_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg322_out;
SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg105_out;
SharedReg198_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg198_out;
SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg737_out;
SharedReg704_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg704_out;
SharedReg706_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg706_out;
SharedReg538_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg538_out;
SharedReg701_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg701_out;
SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg947_out;
SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg737_out;
SharedReg525_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg525_out;
SharedReg1107_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1107_out;
SharedReg314_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg314_out;
SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg105_out;
SharedReg738_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg738_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1108_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg206_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg416_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg322_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg198_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg704_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg706_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg538_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg701_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg947_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg737_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg525_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1107_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg314_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg105_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg738_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg467_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg25_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg703_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg705_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Subtract4_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_2_impl_out,
                 X => Delay1No218_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg211_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg120_out;
SharedReg660_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg660_out;
SharedReg708_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg708_out;
SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg659_out;
SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg659_out;
Delay10No20_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast <= Delay10No20_out;
SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg8_out;
SharedReg422_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg422_out;
SharedReg424_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg424_out;
SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg658_out;
SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg120_out;
SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg707_out;
SharedReg332_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg332_out;
SharedReg116_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg116_out;
SharedReg48_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg48_out;
SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg658_out;
SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg707_out;
SharedReg909_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg909_out;
SharedReg818_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg818_out;
SharedReg743_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg743_out;
SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg707_out;
SharedReg472_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg472_out;
SharedReg809_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg809_out;
SharedReg953_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg953_out;
   MUX_Subtract4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg8_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg422_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg424_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg120_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg332_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg116_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg48_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg658_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg660_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg909_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg818_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg743_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg707_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg472_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg809_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg953_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg708_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg659_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay10No20_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_2_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_0_out,
                 Y => Delay1No218_out);

SharedReg326_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg115_out;
SharedReg708_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg708_out;
SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg955_out;
SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg955_out;
SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg954_out;
SharedReg473_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg473_out;
SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg24_out;
SharedReg709_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg709_out;
SharedReg711_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg711_out;
SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg742_out;
SharedReg219_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg219_out;
SharedReg421_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg421_out;
SharedReg334_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg334_out;
SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg115_out;
SharedReg211_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg211_out;
SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg742_out;
SharedReg710_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg710_out;
SharedReg712_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg712_out;
SharedReg552_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg552_out;
SharedReg707_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg707_out;
SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg954_out;
SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg742_out;
SharedReg539_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg539_out;
SharedReg910_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg910_out;
   MUX_Subtract4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg24_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg709_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg711_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg219_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg421_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg334_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg115_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg211_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg708_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg710_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg712_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg552_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg707_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg742_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg539_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg910_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg955_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg954_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg473_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_2_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Subtract4_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_3_impl_out,
                 X => Delay1No220_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg425_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg425_out;
SharedReg822_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg822_out;
SharedReg747_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg747_out;
SharedReg224_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
SharedReg480_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg480_out;
SharedReg714_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg714_out;
SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg664_out;
SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg664_out;
Delay10No21_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast <= Delay10No21_out;
SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg8_out;
SharedReg427_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg427_out;
SharedReg429_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg429_out;
SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg663_out;
SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg130_out;
SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg713_out;
SharedReg344_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg344_out;
SharedReg126_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg126_out;
SharedReg55_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg55_out;
SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg663_out;
SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg713_out;
SharedReg900_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg900_out;
SharedReg831_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg831_out;
SharedReg748_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg748_out;
SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg713_out;
   MUX_Subtract4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg425_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg822_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg9_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg8_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg427_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg429_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg344_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg747_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg126_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg55_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg663_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg900_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg831_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg748_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg713_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg224_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg480_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg714_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg664_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay10No21_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_3_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_0_out,
                 Y => Delay1No220_out);

SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg713_out;
SharedReg553_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg553_out;
SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg914_out;
SharedReg338_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg338_out;
SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg125_out;
SharedReg714_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg714_out;
SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg915_out;
SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg915_out;
SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg914_out;
SharedReg479_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg479_out;
SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
SharedReg715_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg715_out;
SharedReg717_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg717_out;
SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg747_out;
SharedReg232_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg232_out;
SharedReg426_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg426_out;
SharedReg346_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg346_out;
SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg125_out;
SharedReg224_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg224_out;
SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg747_out;
SharedReg716_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg716_out;
SharedReg718_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg718_out;
SharedReg566_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg566_out;
SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg713_out;
SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg914_out;
   MUX_Subtract4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg553_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg25_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg715_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg717_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg232_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg426_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg346_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg224_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg747_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg716_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg718_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg566_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg713_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg338_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg125_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg714_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg915_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg914_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg479_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_3_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Subtract4_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_4_impl_out,
                 X => Delay1No222_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg844_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg844_out;
SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg720_out;
SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg668_out;
SharedReg900_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg835_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg753_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg753_out;
SharedReg237_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg237_out;
SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg140_out;
SharedReg486_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg486_out;
SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg720_out;
SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg669_out;
SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg669_out;
Delay10No22_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast <= Delay10No22_out;
SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg8_out;
SharedReg432_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg432_out;
SharedReg434_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg434_out;
SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg668_out;
SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg140_out;
SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg719_out;
SharedReg356_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg356_out;
SharedReg136_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg136_out;
SharedReg62_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg62_out;
SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg668_out;
SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg719_out;
SharedReg453_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg453_out;
   MUX_Subtract4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg844_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg669_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay10No22_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg5_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg9_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg8_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg432_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg434_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg356_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg136_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg62_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg668_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg719_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg453_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg900_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg753_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg237_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg140_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg486_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg720_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_4_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_0_out,
                 Y => Delay1No222_out);

SharedReg580_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg580_out;
SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg668_out;
SharedReg754_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg754_out;
SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg668_out;
SharedReg567_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg567_out;
SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg904_out;
SharedReg350_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg350_out;
SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg135_out;
SharedReg720_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg720_out;
SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg905_out;
SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg905_out;
SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg904_out;
SharedReg485_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg485_out;
SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg24_out;
SharedReg721_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg721_out;
SharedReg723_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg723_out;
SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg753_out;
SharedReg245_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg245_out;
SharedReg431_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg431_out;
SharedReg358_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg358_out;
SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg135_out;
SharedReg237_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg237_out;
SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg753_out;
SharedReg722_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg722_out;
SharedReg724_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg724_out;
   MUX_Subtract4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg580_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg485_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg21_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg25_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg24_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg721_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg723_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg754_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg245_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg431_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg358_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg237_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg753_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg722_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg724_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg668_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg567_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg904_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg350_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg135_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg720_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg905_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_4_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Subtract4_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_5_impl_out,
                 X => Delay1No224_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg490_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg490_out;
SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg673_out;
SharedReg456_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg456_out;
SharedReg857_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg857_out;
SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg674_out;
SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg673_out;
SharedReg453_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg453_out;
SharedReg848_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg848_out;
SharedReg932_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg932_out;
SharedReg250_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg250_out;
SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg150_out;
SharedReg492_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg492_out;
SharedReg760_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg760_out;
SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg674_out;
SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg674_out;
Delay10No23_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_16_cast <= Delay10No23_out;
SharedReg1_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg8_out;
SharedReg437_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg437_out;
SharedReg439_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg439_out;
SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg673_out;
SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg150_out;
SharedReg759_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg759_out;
SharedReg368_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg368_out;
SharedReg146_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg146_out;
SharedReg69_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg69_out;
   MUX_Subtract4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg490_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg492_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg760_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay10No23_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg5_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg9_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg8_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg456_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg437_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg439_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg759_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg368_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg146_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg69_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg857_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg674_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg673_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg453_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg848_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg932_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg250_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_5_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_5_impl_0_out,
                 Y => Delay1No224_out);

SharedReg759_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg759_out;
SharedReg762_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg762_out;
SharedReg764_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg764_out;
SharedReg594_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg594_out;
SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg673_out;
SharedReg933_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg673_out;
SharedReg581_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg581_out;
SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg457_out;
SharedReg362_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg362_out;
SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg145_out;
SharedReg760_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg760_out;
SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg458_out;
SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg458_out;
SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg457_out;
SharedReg491_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg491_out;
SharedReg17_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg24_out;
SharedReg761_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg761_out;
SharedReg763_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg763_out;
SharedReg932_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg932_out;
SharedReg258_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg258_out;
SharedReg436_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg436_out;
SharedReg370_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg370_out;
SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg145_out;
SharedReg250_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg250_out;
   MUX_Subtract4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg759_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg762_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg760_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg458_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg491_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg17_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg21_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg25_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg24_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg764_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg761_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg763_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg932_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg258_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg436_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg370_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg145_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg250_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg594_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg673_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg581_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg457_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg362_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_5_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_5_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Subtract4_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_6_impl_out,
                 X => Delay1No226_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg380_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg380_out;
SharedReg156_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
SharedReg76_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg76_out;
SharedReg496_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg496_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg766_out;
SharedReg444_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg444_out;
SharedReg870_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg870_out;
SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg767_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg766_out;
SharedReg440_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg440_out;
SharedReg861_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg861_out;
SharedReg960_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg960_out;
SharedReg263_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg263_out;
SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg160_out;
SharedReg680_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg680_out;
SharedReg921_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg921_out;
SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg767_out;
SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg767_out;
Delay10No24_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_19_cast <= Delay10No24_out;
SharedReg1_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg8_out;
SharedReg498_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg498_out;
SharedReg500_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg500_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg766_out;
SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg160_out;
SharedReg920_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg920_out;
   MUX_Subtract4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg380_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg861_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg960_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg263_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg680_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg921_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay10No24_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg76_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg5_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg9_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg8_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg498_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg500_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg160_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg920_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg496_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg444_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg870_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg767_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg766_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg440_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_6_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_6_impl_0_out,
                 Y => Delay1No226_out);

SharedReg382_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg382_out;
SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg155_out;
SharedReg263_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg766_out;
SharedReg769_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg769_out;
SharedReg771_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg771_out;
SharedReg608_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg608_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg766_out;
SharedReg961_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg961_out;
SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg766_out;
SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg595_out;
SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg445_out;
SharedReg374_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg374_out;
SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg155_out;
SharedReg921_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg921_out;
SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg446_out;
SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg446_out;
SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg445_out;
SharedReg679_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg679_out;
SharedReg17_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg24_out;
SharedReg922_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg922_out;
SharedReg924_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg924_out;
SharedReg960_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg960_out;
SharedReg271_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg271_out;
SharedReg497_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg497_out;
   MUX_Subtract4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg382_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg374_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg155_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg921_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg446_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg445_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg679_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg17_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg263_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg21_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg25_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg24_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg922_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg924_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg960_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg271_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg497_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg769_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg771_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg608_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg961_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg766_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_6_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_6_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Subtract4_7_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Subtract4_7_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Subtract4_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_7_impl_out,
                 X => Delay1No228_out_to_Subtract4_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Subtract4_7_impl_parent_implementedSystem_port_1_cast);

SharedReg683_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg683_out;
SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg772_out;
SharedReg392_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg166_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg166_out;
SharedReg83_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg83_out;
SharedReg642_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg642_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg772_out;
SharedReg637_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg637_out;
SharedReg883_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg883_out;
SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg773_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg772_out;
SharedReg502_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg502_out;
SharedReg874_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg874_out;
SharedReg966_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg966_out;
SharedReg276_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg276_out;
SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg170_out;
SharedReg685_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg685_out;
SharedReg927_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg927_out;
SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg773_out;
SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg773_out;
Delay10No25_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_22_cast <= Delay10No25_out;
SharedReg1_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg8_out;
SharedReg644_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg644_out;
SharedReg646_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg646_out;
   MUX_Subtract4_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg683_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg502_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg874_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg966_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg276_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg170_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg685_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg927_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg773_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay10No25_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg5_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg9_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg8_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg644_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg646_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg392_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg166_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg83_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg642_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg772_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg637_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg883_out_to_MUX_Subtract4_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_7_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_7_impl_0_out,
                 Y => Delay1No228_out);

SharedReg926_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg926_out;
SharedReg284_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg284_out;
SharedReg503_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg503_out;
SharedReg394_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg394_out;
SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg165_out;
SharedReg276_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg276_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg772_out;
SharedReg775_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg775_out;
SharedReg688_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg688_out;
SharedReg622_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg622_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg772_out;
SharedReg967_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg967_out;
SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg772_out;
SharedReg609_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg609_out;
SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg638_out;
SharedReg386_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg386_out;
SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg165_out;
SharedReg927_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg927_out;
SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg639_out;
SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg639_out;
SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg638_out;
SharedReg684_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg684_out;
SharedReg17_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg24_out;
SharedReg928_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg928_out;
SharedReg930_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg930_out;
   MUX_Subtract4_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg926_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg284_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg967_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg609_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg386_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg927_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg639_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg503_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg638_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg684_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg17_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg21_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg25_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg24_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg928_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg930_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg394_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg165_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg276_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg772_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg775_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg688_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg622_out_to_MUX_Subtract4_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_7_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_7_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Subtract4_8_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Subtract4_8_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Subtract4_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_8_impl_out,
                 X => Delay1No230_out_to_Subtract4_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Subtract4_8_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg452_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg452_out;
SharedReg509_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg509_out;
SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg689_out;
SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg180_out;
SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg689_out;
SharedReg404_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg404_out;
SharedReg176_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg90_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg90_out;
SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg689_out;
SharedReg726_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg726_out;
SharedReg972_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg972_out;
SharedReg896_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg896_out;
SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg779_out;
SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg689_out;
SharedReg505_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg505_out;
SharedReg887_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg887_out;
SharedReg778_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg778_out;
SharedReg289_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg289_out;
SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg180_out;
SharedReg728_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg728_out;
SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg727_out;
SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg779_out;
SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg727_out;
Delay10No26_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_26_cast <= Delay10No26_out;
SharedReg1_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg5_out;
   MUX_Subtract4_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg726_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg972_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg896_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg505_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg887_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg778_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg289_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg452_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg728_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg779_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg727_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay10No26_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg5_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg509_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg180_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg689_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg404_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg90_out_to_MUX_Subtract4_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_8_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_8_impl_0_out,
                 Y => Delay1No230_out);

SharedReg25_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg24_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg728_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg728_out;
SharedReg782_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg782_out;
SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg778_out;
SharedReg297_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
SharedReg451_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg451_out;
SharedReg406_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg406_out;
SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg175_out;
SharedReg289_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg289_out;
SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg778_out;
SharedReg729_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg729_out;
SharedReg731_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg731_out;
SharedReg636_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg636_out;
SharedReg726_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg726_out;
SharedReg973_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg973_out;
SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg778_out;
SharedReg623_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg623_out;
SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg980_out;
SharedReg398_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg398_out;
SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg175_out;
SharedReg779_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg779_out;
SharedReg981_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg981_out;
SharedReg974_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg974_out;
SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg980_out;
SharedReg690_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg690_out;
SharedReg17_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg17_out;
SharedReg21_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg21_out;
   MUX_Subtract4_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg729_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg731_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg636_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg726_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg973_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg623_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg398_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg728_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg779_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg981_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg974_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg980_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg690_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg17_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg21_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg782_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg778_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg297_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg451_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg406_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg175_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg289_out_to_MUX_Subtract4_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract4_8_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_8_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product34_4_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product34_4_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product34_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product34_4_impl_out,
                 X => Delay1No232_out_to_Product34_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product34_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1200_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1229_out;
SharedReg1203_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1204_out;
SharedReg238_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg1206_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1206_out;
SharedReg62_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg62_out;
SharedReg1207_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1207_out;
SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1134_out;
SharedReg1137_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1275_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1259_out;
SharedReg1136_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1136_out;
SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1134_out;
SharedReg1183_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1288_out;
SharedReg1185_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1185_out;
SharedReg341_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg341_out;
SharedReg1187_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1218_out;
SharedReg570_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg570_out;
SharedReg1268_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1268_out;
SharedReg1278_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1278_out;
SharedReg1252_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1252_out;
   MUX_Product34_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1200_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1201_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1275_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1281_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1259_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1136_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1183_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1288_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1185_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg341_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1229_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1187_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1188_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1189_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1218_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg570_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1268_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1278_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1252_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1203_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1204_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg238_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1206_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg62_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1207_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1134_out_to_MUX_Product34_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product34_4_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_4_impl_0_out,
                 Y => Delay1No232_out);

SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg238_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg135_out;
SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg61_out;
SharedReg1232_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1232_out;
SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg61_out;
SharedReg1234_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1234_out;
SharedReg60_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
SharedReg1245_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1280_out;
SharedReg1138_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1138_out;
SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1136_out;
SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1136_out;
SharedReg1260_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1287_out;
SharedReg224_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg224_out;
SharedReg1026_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1026_out;
SharedReg825_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg825_out;
SharedReg1214_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1214_out;
SharedReg558_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg558_out;
SharedReg341_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg341_out;
SharedReg343_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg343_out;
SharedReg58_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg58_out;
SharedReg1248_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1248_out;
SharedReg1147_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1147_out;
SharedReg1042_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1042_out;
SharedReg1046_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1046_out;
   MUX_Product34_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1280_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1138_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1136_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1260_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1287_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg224_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1026_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg825_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1214_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg558_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg341_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg343_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg58_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1248_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1147_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1042_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1046_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg135_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1232_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg61_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1234_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1245_out_to_MUX_Product34_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product34_4_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_4_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product34_5_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product34_5_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product34_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product34_5_impl_out,
                 X => Delay1No234_out_to_Product34_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product34_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1142_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1142_out;
SharedReg1263_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1272_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg837_out;
SharedReg1144_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1144_out;
SharedReg1202_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1202_out;
SharedReg1145_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1145_out;
SharedReg1149_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1149_out;
SharedReg1205_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1205_out;
SharedReg1037_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1037_out;
SharedReg1279_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1245_out;
SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg837_out;
SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg837_out;
SharedReg1276_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1286_out;
SharedReg135_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg135_out;
SharedReg1212_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1212_out;
SharedReg239_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg239_out;
SharedReg1214_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1214_out;
SharedReg138_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg138_out;
SharedReg1188_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1218_out;
SharedReg584_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg584_out;
   MUX_Product34_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1142_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1279_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1244_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1245_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1276_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1250_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1251_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1286_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg135_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1212_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg239_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1214_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg138_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1188_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1189_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1218_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg584_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg837_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1144_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1202_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1145_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1149_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1205_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1037_out_to_MUX_Product34_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product34_5_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_5_impl_0_out,
                 Y => Delay1No234_out);

SharedReg1262_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1262_out;
SharedReg1038_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1038_out;
SharedReg1056_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1056_out;
SharedReg1265_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1231_out;
SharedReg68_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg68_out;
SharedReg1233_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1237_out;
SharedReg251_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg251_out;
SharedReg1219_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1219_out;
SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1037_out;
SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1037_out;
SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1037_out;
SharedReg1280_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1223_out;
SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1144_out;
SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1144_out;
SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1144_out;
SharedReg1142_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1142_out;
SharedReg1211_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1211_out;
SharedReg61_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg61_out;
SharedReg1213_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1213_out;
SharedReg351_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg351_out;
SharedReg1215_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1215_out;
SharedReg353_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg353_out;
SharedReg355_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg355_out;
SharedReg65_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg65_out;
SharedReg1248_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1248_out;
   MUX_Product34_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1262_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1038_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1037_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1280_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1223_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1144_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1142_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1211_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1056_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg61_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1213_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg351_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1215_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg353_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg355_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg65_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1248_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1265_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1231_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg68_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1233_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1237_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg251_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1219_out_to_MUX_Product34_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product34_5_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_5_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product10_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_3_impl_out,
                 X => Delay1No236_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1203_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1204_out;
SharedReg225_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg225_out;
SharedReg1206_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1206_out;
SharedReg55_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg55_out;
SharedReg1207_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1207_out;
SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1126_out;
SharedReg1129_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1129_out;
SharedReg1275_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1259_out;
SharedReg1128_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1128_out;
SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1126_out;
SharedReg1183_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1288_out;
SharedReg1185_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1185_out;
SharedReg329_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg329_out;
SharedReg1187_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1218_out;
SharedReg1236_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1236_out;
SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1126_out;
SharedReg1263_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1263_out;
SharedReg1272_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1272_out;
SharedReg1200_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1200_out;
SharedReg1201_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1201_out;
SharedReg1229_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1229_out;
   MUX_Product10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1203_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1204_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1259_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1128_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1183_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1288_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1185_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg329_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1187_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1188_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1189_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg225_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1218_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1236_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1263_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1272_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1200_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1201_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1229_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1206_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg55_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1207_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1126_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1129_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1275_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1281_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product10_3_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_3_impl_0_out,
                 Y => Delay1No236_out);

SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg54_out;
SharedReg1232_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1232_out;
SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg54_out;
SharedReg1234_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1234_out;
SharedReg53_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg53_out;
SharedReg1245_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1280_out;
SharedReg1130_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1130_out;
SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1128_out;
SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1128_out;
SharedReg1260_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1287_out;
SharedReg211_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg211_out;
SharedReg1013_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1013_out;
SharedReg812_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg812_out;
SharedReg1214_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1214_out;
SharedReg544_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg544_out;
SharedReg329_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg329_out;
SharedReg331_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg331_out;
SharedReg51_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg51_out;
SharedReg52_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg52_out;
SharedReg1262_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1262_out;
SharedReg1012_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1012_out;
SharedReg1030_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1030_out;
SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg125_out;
SharedReg225_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg225_out;
SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg54_out;
   MUX_Product10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1260_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1287_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg211_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1013_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg812_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1214_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg544_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg329_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg331_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1232_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg51_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg52_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1262_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1012_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1030_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg125_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg225_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg54_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1234_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg53_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1245_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1280_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1130_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1128_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product10_3_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_3_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Product10_4_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Product10_4_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Product10_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_4_impl_out,
                 X => Delay1No238_out_to_Product10_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Product10_4_impl_parent_implementedSystem_port_1_cast);

SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg824_out;
SharedReg1136_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1136_out;
SharedReg1202_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1202_out;
SharedReg1137_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1141_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1141_out;
SharedReg1205_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1205_out;
SharedReg1024_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1024_out;
SharedReg1279_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1245_out;
SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg824_out;
SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg824_out;
SharedReg1276_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1286_out;
SharedReg125_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg125_out;
SharedReg1212_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1212_out;
SharedReg226_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg226_out;
SharedReg1214_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1214_out;
SharedReg128_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg1216_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1216_out;
SharedReg342_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg342_out;
SharedReg1190_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1190_out;
SharedReg1236_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1236_out;
SharedReg1134_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1134_out;
SharedReg1263_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1263_out;
SharedReg1272_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1272_out;
   MUX_Product10_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1136_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1276_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1250_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1251_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1286_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg125_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1212_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg226_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1214_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1202_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1216_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg342_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1190_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1236_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1134_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1263_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1272_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1141_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1205_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1024_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1279_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1244_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1245_out_to_MUX_Product10_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product10_4_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_4_impl_0_out,
                 Y => Delay1No238_out);

SharedReg1265_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1231_out;
SharedReg61_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg1233_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1237_out;
SharedReg238_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg1219_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1219_out;
SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1024_out;
SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1024_out;
SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1024_out;
SharedReg1280_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1223_out;
SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1136_out;
SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1136_out;
SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1136_out;
SharedReg1134_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1134_out;
SharedReg1211_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1211_out;
SharedReg54_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg54_out;
SharedReg1213_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1213_out;
SharedReg339_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg339_out;
SharedReg1215_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1215_out;
SharedReg57_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg57_out;
SharedReg1217_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1217_out;
SharedReg58_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg58_out;
SharedReg59_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg59_out;
SharedReg1262_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1262_out;
SharedReg1025_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1025_out;
SharedReg1043_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1043_out;
   MUX_Product10_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1265_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1231_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1280_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1223_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1136_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1134_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1211_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg54_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1213_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg339_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1215_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg57_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1217_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg58_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg59_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1262_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1025_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1043_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1233_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1237_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg238_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1219_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1024_out_to_MUX_Product10_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product10_4_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_4_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Product28_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_6_impl_out,
                 X => Delay1No240_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1285_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1187_out;
SharedReg1216_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1216_out;
SharedReg1189_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1208_out;
SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg374_out;
SharedReg1201_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1255_out;
SharedReg1160_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1160_out;
SharedReg1257_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1235_out;
SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg155_out;
SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg155_out;
SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg374_out;
SharedReg1242_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1196_out;
SharedReg1224_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1225_out;
SharedReg1199_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1184_out;
SharedReg265_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg265_out;
   MUX_Product28_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1285_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1187_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1257_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1205_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1206_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1209_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1235_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1242_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1216_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1196_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1224_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1225_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1199_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1286_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1183_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1184_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg265_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1189_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1218_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1208_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg374_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1201_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1255_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1160_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_6_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_6_impl_0_out,
                 Y => Delay1No240_out);

SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1159_out;
SharedReg158_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg158_out;
SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg378_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg378_out;
SharedReg268_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg268_out;
SharedReg80_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg80_out;
SharedReg1227_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1227_out;
SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg75_out;
SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg863_out;
SharedReg1265_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1265_out;
SharedReg1065_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1065_out;
SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1161_out;
SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1161_out;
SharedReg1165_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1165_out;
SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1159_out;
SharedReg1219_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1222_out;
SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1159_out;
SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg863_out;
SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg78_out;
SharedReg157_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg157_out;
SharedReg76_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg76_out;
SharedReg1063_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1063_out;
SharedReg155_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg155_out;
SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg75_out;
SharedReg1213_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1213_out;
   MUX_Product28_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1065_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1161_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1165_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1219_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1220_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1221_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1222_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1159_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg78_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg157_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg76_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1063_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg155_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1213_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg378_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg268_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg80_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1227_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg75_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg863_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1265_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_6_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_6_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product28_7_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product28_7_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product28_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_7_impl_out,
                 X => Delay1No242_out_to_Product28_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product28_7_impl_parent_implementedSystem_port_1_cast);

SharedReg1183_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1184_out;
SharedReg278_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg278_out;
SharedReg1285_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1285_out;
SharedReg1187_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1187_out;
SharedReg1216_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1216_out;
SharedReg1189_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1208_out;
SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg386_out;
SharedReg1201_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1201_out;
SharedReg1255_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1255_out;
SharedReg1168_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1168_out;
SharedReg1257_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1257_out;
SharedReg1205_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1206_out;
SharedReg1209_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1209_out;
SharedReg1235_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1235_out;
SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg165_out;
SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg165_out;
SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg386_out;
SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg386_out;
SharedReg1242_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1242_out;
SharedReg1196_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1196_out;
SharedReg169_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg169_out;
SharedReg83_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg83_out;
SharedReg1199_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1286_out;
   MUX_Product28_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1183_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1184_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1201_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1255_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1168_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1257_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1205_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1206_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1209_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1235_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg165_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg278_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1242_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1196_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg169_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg83_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1199_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1286_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1285_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1187_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1216_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1189_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1218_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1208_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg386_out_to_MUX_Product28_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_7_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_7_impl_0_out,
                 Y => Delay1No242_out);

SharedReg165_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg1213_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1213_out;
SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1167_out;
SharedReg168_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg168_out;
SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg85_out;
SharedReg390_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg390_out;
SharedReg281_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg281_out;
SharedReg87_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg87_out;
SharedReg1227_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1227_out;
SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg82_out;
SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg876_out;
SharedReg1265_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1265_out;
SharedReg1078_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1078_out;
SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1169_out;
SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1169_out;
SharedReg1173_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1173_out;
SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1167_out;
SharedReg1219_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1219_out;
SharedReg1220_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1220_out;
SharedReg1221_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1221_out;
SharedReg1222_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1222_out;
SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1167_out;
SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg876_out;
SharedReg1224_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1225_out;
SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg85_out;
SharedReg1166_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1166_out;
   MUX_Product28_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg82_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1265_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1078_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1169_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1173_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1219_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1220_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1213_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1221_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1222_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg876_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1224_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1225_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1166_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1167_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg168_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg85_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg390_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg281_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg87_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1227_out_to_MUX_Product28_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product28_7_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_7_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product42_5_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product42_5_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product42_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_5_impl_out,
                 X => Delay1No244_out_to_Product42_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product42_5_impl_parent_implementedSystem_port_1_cast);

SharedReg366_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg366_out;
SharedReg1190_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1190_out;
SharedReg1236_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1236_out;
SharedReg1253_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1254_out;
SharedReg850_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg850_out;
SharedReg1256_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1237_out;
SharedReg1054_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1054_out;
SharedReg1191_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1223_out;
SharedReg149_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg149_out;
SharedReg69_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg69_out;
SharedReg1199_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1286_out;
SharedReg1183_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1183_out;
SharedReg1184_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1184_out;
SharedReg252_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg252_out;
SharedReg1214_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1214_out;
SharedReg148_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg148_out;
SharedReg1188_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1188_out;
   MUX_Product42_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg366_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1190_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1237_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1054_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1191_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1273_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1240_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1241_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1274_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1223_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg149_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg69_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1236_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1199_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1286_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1183_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1184_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg252_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1214_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg148_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1188_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1253_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1254_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg850_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1232_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1233_out_to_MUX_Product42_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product42_5_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_5_impl_0_out,
                 Y => Delay1No244_out);

SharedReg1217_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1217_out;
SharedReg72_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg73_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg73_out;
SharedReg1150_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1150_out;
SharedReg1051_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1051_out;
SharedReg1264_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1264_out;
SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg850_out;
SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1052_out;
SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1052_out;
SharedReg1152_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1152_out;
SharedReg1062_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1062_out;
SharedReg1235_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1235_out;
SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1050_out;
SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1050_out;
SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1050_out;
SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1050_out;
SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg850_out;
SharedReg583_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg583_out;
SharedReg1224_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1225_out;
SharedReg71_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg71_out;
SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1050_out;
SharedReg145_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg145_out;
SharedReg68_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg68_out;
SharedReg1213_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1213_out;
SharedReg363_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg363_out;
SharedReg1215_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1215_out;
SharedReg365_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg365_out;
   MUX_Product42_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1217_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1062_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1235_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg583_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1224_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1225_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg73_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg71_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1050_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg145_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg68_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1213_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg363_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1215_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg365_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1150_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1051_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1264_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg850_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1052_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1152_out_to_MUX_Product42_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product42_5_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_5_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product213_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_0_impl_out,
                 X => Delay1No246_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1245_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1245_out;
SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg785_out;
SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg785_out;
SharedReg1276_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1286_out;
SharedReg95_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg95_out;
SharedReg1212_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1212_out;
SharedReg187_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg187_out;
SharedReg1214_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1214_out;
SharedReg98_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg98_out;
SharedReg1216_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1216_out;
SharedReg306_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg306_out;
SharedReg1190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1190_out;
SharedReg1208_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1208_out;
SharedReg1253_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1266_out;
SharedReg1205_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1237_out;
SharedReg989_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg989_out;
SharedReg985_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg985_out;
SharedReg1279_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1244_out;
   MUX_Product213_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1245_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1214_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1216_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg306_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1190_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1208_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1253_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1254_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1255_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1256_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg785_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1266_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1205_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1233_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1237_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg989_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg985_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1279_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1244_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1276_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1250_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1251_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1286_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg95_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1212_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg187_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_0_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_0_out,
                 Y => Delay1No246_out);

SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg985_out;
SharedReg1280_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1223_out;
SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1112_out;
SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg1211_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1211_out;
SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg1213_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1213_out;
SharedReg303_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg303_out;
SharedReg1215_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1215_out;
SharedReg36_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg36_out;
SharedReg1217_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1217_out;
SharedReg37_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg37_out;
SharedReg38_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg38_out;
SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1110_out;
SharedReg986_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg986_out;
SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg785_out;
SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg785_out;
SharedReg987_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg987_out;
SharedReg1113_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1113_out;
SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1112_out;
SharedReg997_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg997_out;
SharedReg1235_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1235_out;
SharedReg1219_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1219_out;
SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg985_out;
SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg985_out;
   MUX_Product213_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1280_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg303_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1215_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg36_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1217_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg37_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg38_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg986_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg785_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1223_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg987_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1113_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg997_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1235_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1219_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg985_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1211_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1213_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_0_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product213_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_1_impl_out,
                 X => Delay1No248_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast);

SharedReg998_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg998_out;
SharedReg1279_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1245_out;
SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg798_out;
SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg798_out;
SharedReg1276_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1286_out;
SharedReg105_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg105_out;
SharedReg1212_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1212_out;
SharedReg200_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg200_out;
SharedReg1214_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1214_out;
SharedReg108_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg108_out;
SharedReg1216_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1216_out;
SharedReg318_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg318_out;
SharedReg1190_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1190_out;
SharedReg1208_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1208_out;
SharedReg1253_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1254_out;
SharedReg1255_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1232_out;
SharedReg1121_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1121_out;
SharedReg1125_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1125_out;
SharedReg1205_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1205_out;
   MUX_Product213_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg998_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1279_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg105_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1212_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg200_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1214_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg108_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1216_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg318_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1190_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1208_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1253_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1244_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1254_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1255_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1256_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1266_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1232_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1121_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1125_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1205_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1245_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg798_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1276_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1250_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1251_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1286_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_1_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_1_impl_0_out,
                 Y => Delay1No248_out);

SharedReg1219_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1219_out;
SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg998_out;
SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg998_out;
SharedReg1280_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1223_out;
SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1120_out;
SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1120_out;
SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg1211_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1211_out;
SharedReg40_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg40_out;
SharedReg1213_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1213_out;
SharedReg315_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg315_out;
SharedReg1215_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1215_out;
SharedReg43_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg43_out;
SharedReg1217_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1217_out;
SharedReg44_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg44_out;
SharedReg45_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg45_out;
SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1118_out;
SharedReg999_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg999_out;
SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg798_out;
SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg798_out;
SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1000_out;
SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1000_out;
SharedReg1233_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1237_out;
SharedReg212_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg212_out;
   MUX_Product213_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1219_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1211_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg40_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1213_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg315_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1215_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg43_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1217_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg44_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg45_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg999_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg798_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1000_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1233_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1237_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg212_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg998_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1280_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1223_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1120_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_1_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_1_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Product213_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_2_impl_out,
                 X => Delay1No250_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1129_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1133_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1133_out;
SharedReg1205_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1205_out;
SharedReg1011_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1011_out;
SharedReg1279_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1279_out;
SharedReg1244_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1245_out;
SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg811_out;
SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg811_out;
SharedReg1276_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1251_out;
SharedReg1286_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1286_out;
SharedReg115_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg115_out;
SharedReg1212_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1212_out;
SharedReg213_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg213_out;
SharedReg1214_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1214_out;
SharedReg118_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg118_out;
SharedReg1216_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1216_out;
SharedReg330_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg330_out;
SharedReg1190_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1190_out;
SharedReg1208_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1208_out;
SharedReg1253_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1254_out;
SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg811_out;
SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg811_out;
SharedReg1128_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1128_out;
SharedReg1202_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1202_out;
   MUX_Product213_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1133_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1250_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1251_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1286_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg115_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1212_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg213_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1214_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg118_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1216_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg330_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1205_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1190_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1208_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1253_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1254_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1128_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1202_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1011_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1279_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1244_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1245_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg811_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1276_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_2_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_2_impl_0_out,
                 Y => Delay1No250_out);

SharedReg1233_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1237_out;
SharedReg225_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg225_out;
SharedReg1219_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1219_out;
SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1011_out;
SharedReg1280_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1280_out;
SharedReg1223_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1223_out;
SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1128_out;
SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1128_out;
SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1128_out;
SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1126_out;
SharedReg1211_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1211_out;
SharedReg47_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg47_out;
SharedReg1213_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1213_out;
SharedReg327_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg327_out;
SharedReg1215_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1215_out;
SharedReg50_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg50_out;
SharedReg1217_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1217_out;
SharedReg51_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg51_out;
SharedReg52_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg52_out;
SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1126_out;
SharedReg1012_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1012_out;
SharedReg1264_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1231_out;
SharedReg54_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg54_out;
   MUX_Product213_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1233_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1237_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1211_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg47_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1213_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg327_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1215_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg50_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1217_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg225_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg51_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg52_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1126_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1012_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1264_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1265_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1231_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg54_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1219_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1011_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1280_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1223_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1128_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_2_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_2_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Product213_6_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Product213_6_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Product213_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_6_impl_out,
                 X => Delay1No252_out_to_Product213_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Product213_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1214_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1214_out;
SharedReg158_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg158_out;
SharedReg1188_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1188_out;
SharedReg378_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg378_out;
SharedReg1190_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1190_out;
SharedReg1236_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1236_out;
SharedReg1253_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1254_out;
SharedReg863_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg863_out;
SharedReg1256_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1237_out;
SharedReg1067_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1067_out;
SharedReg1191_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1223_out;
SharedReg159_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg159_out;
SharedReg76_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg76_out;
SharedReg1199_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1199_out;
SharedReg1286_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1286_out;
SharedReg155_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg155_out;
SharedReg1212_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1212_out;
SharedReg1185_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1185_out;
   MUX_Product213_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1214_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1266_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1232_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1233_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1237_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1067_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1191_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1273_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1240_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1241_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1274_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1188_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1223_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg159_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg76_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1199_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1286_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg155_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1212_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1185_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg378_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1190_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1236_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1253_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1254_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg863_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1256_out_to_MUX_Product213_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_6_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_6_impl_0_out,
                 Y => Delay1No252_out);

SharedReg375_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg375_out;
SharedReg1215_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1215_out;
SharedReg377_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg1217_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1217_out;
SharedReg79_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg79_out;
SharedReg80_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg80_out;
SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1064_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1064_out;
SharedReg1264_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg863_out;
SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1065_out;
SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1065_out;
SharedReg1160_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1160_out;
SharedReg1075_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1075_out;
SharedReg1235_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1235_out;
SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1063_out;
SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1063_out;
SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1063_out;
SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1063_out;
SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg863_out;
SharedReg597_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg597_out;
SharedReg1224_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1224_out;
SharedReg1225_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1225_out;
SharedReg78_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg78_out;
SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1158_out;
SharedReg1211_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1211_out;
SharedReg75_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg75_out;
SharedReg864_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg864_out;
   MUX_Product213_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg375_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1215_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1065_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1160_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1075_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1235_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1063_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg377_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg597_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1224_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1225_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg78_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1211_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg75_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg864_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1217_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg79_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg80_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1064_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg863_out_to_MUX_Product213_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_6_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_6_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product213_7_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product213_7_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product213_7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_7_impl_out,
                 X => Delay1No254_out_to_Product213_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product213_7_impl_parent_implementedSystem_port_1_cast);

SharedReg165_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg1212_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1212_out;
SharedReg1185_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1185_out;
SharedReg1214_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1214_out;
SharedReg168_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg168_out;
SharedReg1188_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1188_out;
SharedReg390_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg390_out;
SharedReg1190_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1190_out;
SharedReg1236_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1236_out;
SharedReg1253_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1253_out;
SharedReg1254_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1254_out;
SharedReg876_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg876_out;
SharedReg1256_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1266_out;
SharedReg1232_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1232_out;
SharedReg1233_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1237_out;
SharedReg1080_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1080_out;
SharedReg1191_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1273_out;
SharedReg1240_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1240_out;
SharedReg1241_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1241_out;
SharedReg1274_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1274_out;
SharedReg1223_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1223_out;
SharedReg1276_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1250_out;
SharedReg1251_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1251_out;
SharedReg1166_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1166_out;
   MUX_Product213_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1212_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1254_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg876_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1266_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1232_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1233_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1237_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1080_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1191_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1273_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1185_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1240_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1241_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1274_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1223_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1276_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1250_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1251_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1166_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1214_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg168_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1188_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg390_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1190_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1236_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1253_out_to_MUX_Product213_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_7_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_7_impl_0_out,
                 Y => Delay1No254_out);

SharedReg1211_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1211_out;
SharedReg82_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg877_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg877_out;
SharedReg387_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
SharedReg1215_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1215_out;
SharedReg389_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg389_out;
SharedReg1217_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1217_out;
SharedReg86_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg86_out;
SharedReg87_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg87_out;
SharedReg1166_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1166_out;
SharedReg1077_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1077_out;
SharedReg1264_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1264_out;
SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg876_out;
SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1078_out;
SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1078_out;
SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1168_out;
SharedReg1088_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1088_out;
SharedReg1235_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1235_out;
SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1076_out;
SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1076_out;
SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1076_out;
SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1076_out;
SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg876_out;
SharedReg611_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg611_out;
SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1168_out;
SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1168_out;
SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1168_out;
SharedReg1287_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1287_out;
   MUX_Product213_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1211_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1077_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1264_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1078_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1088_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1235_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg877_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1076_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg876_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg611_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1168_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1287_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg387_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1215_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg389_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1217_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg86_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg87_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1166_out_to_MUX_Product213_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product213_7_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_7_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product313_8_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product313_8_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product313_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_8_impl_out,
                 X => Delay1No256_out_to_Product313_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product313_8_impl_parent_implementedSystem_port_1_cast);

SharedReg1276_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1276_out;
SharedReg1250_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1250_out;
SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1176_out;
SharedReg1286_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1286_out;
SharedReg175_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg1288_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1288_out;
SharedReg291_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg291_out;
SharedReg1214_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1214_out;
SharedReg1187_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1187_out;
SharedReg1216_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1216_out;
SharedReg402_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg402_out;
SharedReg1218_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1218_out;
SharedReg1208_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1208_out;
SharedReg1253_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1253_out;
SharedReg1263_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1263_out;
SharedReg1255_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1255_out;
SharedReg1256_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1256_out;
SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1176_out;
SharedReg1205_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1205_out;
SharedReg1233_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1237_out;
SharedReg1235_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1235_out;
SharedReg1191_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1191_out;
SharedReg1273_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1273_out;
SharedReg1244_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1244_out;
SharedReg1245_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1245_out;
SharedReg889_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg889_out;
SharedReg1275_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1275_out;
   MUX_Product313_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1276_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1250_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg402_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1218_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1208_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1253_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1263_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1255_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1256_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1205_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1233_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1176_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1237_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1235_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1191_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1273_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1244_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1245_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg889_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1275_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1286_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1288_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg291_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1214_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1187_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1216_out_to_MUX_Product313_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product313_8_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_8_impl_0_out,
                 Y => Delay1No256_out);

SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1176_out;
SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1176_out;
SharedReg1260_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1260_out;
SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1174_out;
SharedReg1211_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1211_out;
SharedReg1091_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1091_out;
SharedReg1213_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1213_out;
SharedReg399_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg399_out;
SharedReg628_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg628_out;
SharedReg92_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg92_out;
SharedReg1217_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1217_out;
SharedReg93_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg93_out;
SharedReg94_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg94_out;
SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1174_out;
SharedReg1090_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1090_out;
SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg889_out;
SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg889_out;
SharedReg1231_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1231_out;
SharedReg1177_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1177_out;
SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1176_out;
SharedReg1101_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1101_out;
SharedReg1175_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1175_out;
SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1089_out;
SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1089_out;
SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1089_out;
SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1089_out;
SharedReg1280_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1280_out;
SharedReg1178_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1178_out;
   MUX_Product313_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1217_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg93_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg94_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1090_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg889_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1231_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1177_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1176_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1260_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1101_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1175_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1089_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1280_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1178_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1174_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1211_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1091_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1213_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg399_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg628_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg92_out_to_MUX_Product313_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product313_8_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_8_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product316_8_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product316_8_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product316_8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product316_8_impl_out,
                 X => Delay1No258_out_to_Product316_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product316_8_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg1181_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1181_out;
SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1174_out;
SharedReg1089_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1089_out;
SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1177_out;
SharedReg1093_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1093_out;
SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg889_out;
SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg889_out;
SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1177_out;
SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1174_out;
SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1174_out;
SharedReg1281_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1281_out;
SharedReg1279_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1279_out;
SharedReg1259_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1259_out;
SharedReg1236_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1236_out;
SharedReg1232_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1232_out;
SharedReg1183_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1183_out;
SharedReg1188_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1189_out;
SharedReg1185_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1185_out;
   MUX_Product316_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_20_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1181_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1281_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1279_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1259_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1236_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1232_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1183_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1188_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1189_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1185_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1089_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1093_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg889_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1177_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1174_out_to_MUX_Product316_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product316_8_impl_0_LUT_out,
                 oMux => MUX_Product316_8_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_8_impl_0_out,
                 Y => Delay1No258_out);

SharedReg94_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg403_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg289_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg289_out;
SharedReg401_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg401_out;
SharedReg890_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg890_out;
SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1176_out;
SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1176_out;
SharedReg1089_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1089_out;
SharedReg1091_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1091_out;
SharedReg1219_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1219_out;
SharedReg1245_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1280_out;
SharedReg1265_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1265_out;
SharedReg1237_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1237_out;
SharedReg1235_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1235_out;
SharedReg1264_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1264_out;
SharedReg1262_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1262_out;
SharedReg1233_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1233_out;
SharedReg1214_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1214_out;
SharedReg1287_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1287_out;
   MUX_Product316_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_20_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1245_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1280_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1265_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1237_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1235_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1264_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1262_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1233_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1214_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1287_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg289_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg890_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1176_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1089_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1091_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1219_out_to_MUX_Product316_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product316_8_impl_1_LUT_out,
                 oMux => MUX_Product316_8_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_8_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Subtract18_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_0_impl_out,
                 X => Delay1No260_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg696_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg696_out;
SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg734_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg734_out;
SharedReg648_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg648_out;
SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg939_out;
SharedReg788_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg788_out;
SharedReg940_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg940_out;
SharedReg789_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg789_out;
SharedReg986_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg986_out;
SharedReg1112_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1112_out;
SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg514_out;
SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg514_out;
SharedReg98_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg98_out;
SharedReg194_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg194_out;
SharedReg994_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg994_out;
SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg939_out;
SharedReg522_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg522_out;
SharedReg304_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg304_out;
SharedReg511_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg511_out;
SharedReg518_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg518_out;
SharedReg515_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg515_out;
SharedReg651_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg651_out;
SharedReg192_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg192_out;
SharedReg520_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg520_out;
SharedReg996_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg996_out;
   MUX_Subtract18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg696_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg789_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg986_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1112_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg514_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg98_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg194_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg994_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg522_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg13_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg304_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg511_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg518_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg515_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg651_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg192_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg520_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg996_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg10_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg648_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg939_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg788_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg940_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_0_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_0_impl_0_out,
                 Y => Delay1No260_out);

SharedReg1103_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1103_out;
SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg460_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg460_out;
SharedReg939_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg939_out;
SharedReg941_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg941_out;
SharedReg992_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg992_out;
SharedReg1102_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1102_out;
SharedReg793_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg793_out;
SharedReg1110_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
SharedReg985_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg985_out;
SharedReg784_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg784_out;
SharedReg512_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg512_out;
SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg302_out;
Delay44No_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_17_cast <= Delay44No_out;
Delay45No18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_18_cast <= Delay45No18_out;
SharedReg944_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg944_out;
SharedReg523_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg523_out;
SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg302_out;
SharedReg785_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg785_out;
SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg511_out;
SharedReg783_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg783_out;
SharedReg1104_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1104_out;
SharedReg304_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg304_out;
SharedReg988_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg988_out;
SharedReg786_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg786_out;
   MUX_Subtract18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1103_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg793_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg985_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg784_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg512_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay44No_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay45No18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg944_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg523_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg29_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg302_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg785_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg783_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1104_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg304_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg988_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg786_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg26_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg460_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg939_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg941_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg992_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1102_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_0_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_0_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Subtract18_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_1_impl_out,
                 X => Delay1No262_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg205_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg205_out;
SharedReg534_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg1009_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1009_out;
SharedReg654_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg654_out;
SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg739_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg739_out;
SharedReg653_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg653_out;
SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg946_out;
SharedReg801_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg947_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg947_out;
SharedReg802_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg802_out;
SharedReg999_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg999_out;
SharedReg1120_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1120_out;
SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg528_out;
SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg528_out;
SharedReg108_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg108_out;
SharedReg207_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg207_out;
SharedReg1007_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1007_out;
SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg946_out;
SharedReg536_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg536_out;
SharedReg316_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg316_out;
SharedReg525_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg525_out;
SharedReg532_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg532_out;
SharedReg529_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg529_out;
SharedReg656_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg656_out;
   MUX_Subtract18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg205_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg947_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg802_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg999_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1120_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg528_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg108_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg207_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1009_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1007_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg946_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg536_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg316_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg525_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg532_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg529_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg656_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg654_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg10_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg739_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg653_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_1_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_1_impl_0_out,
                 Y => Delay1No262_out);

SharedReg316_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg316_out;
SharedReg1001_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg799_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg799_out;
SharedReg947_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg947_out;
SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg466_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg466_out;
SharedReg946_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg946_out;
SharedReg948_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg948_out;
SharedReg1005_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1005_out;
SharedReg1106_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1106_out;
SharedReg806_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg806_out;
SharedReg1118_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1118_out;
SharedReg998_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg998_out;
SharedReg797_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg797_out;
SharedReg526_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg526_out;
SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg314_out;
Delay44No1_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_20_cast <= Delay44No1_out;
Delay45No19_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_21_cast <= Delay45No19_out;
SharedReg951_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg951_out;
SharedReg537_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg537_out;
SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg314_out;
SharedReg798_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg798_out;
SharedReg525_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg525_out;
SharedReg796_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg796_out;
SharedReg1108_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1108_out;
   MUX_Subtract18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg316_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg948_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1005_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1106_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg806_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1118_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg998_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg797_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg526_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay44No1_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg799_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay45No19_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg951_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg537_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg314_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg798_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg525_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg796_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1108_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg947_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg26_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg466_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg946_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_1_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_1_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Subtract18_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_2_impl_out,
                 X => Delay1No264_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg546_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg546_out;
SharedReg543_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg543_out;
SharedReg661_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg661_out;
SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg548_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg1022_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1022_out;
SharedReg659_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg659_out;
SharedReg2_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg12_out;
SharedReg744_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg744_out;
SharedReg658_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg658_out;
SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg953_out;
SharedReg814_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg814_out;
SharedReg954_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg954_out;
SharedReg815_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg815_out;
SharedReg1012_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1012_out;
SharedReg1128_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1128_out;
SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg542_out;
SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg542_out;
SharedReg118_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg118_out;
SharedReg220_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg220_out;
SharedReg1020_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1020_out;
SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg953_out;
SharedReg550_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg550_out;
SharedReg328_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg328_out;
SharedReg539_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg539_out;
   MUX_Subtract18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg546_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg543_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg12_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg744_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg658_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg814_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg954_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg815_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1012_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1128_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg661_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg542_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg118_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg220_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1020_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg953_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg550_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg328_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg539_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1022_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg659_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg2_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg10_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_2_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_2_impl_0_out,
                 Y => Delay1No264_out);

SharedReg539_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg539_out;
SharedReg809_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg809_out;
SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg955_out;
SharedReg328_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg1014_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1014_out;
SharedReg812_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg812_out;
SharedReg954_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg954_out;
SharedReg18_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg28_out;
SharedReg472_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg472_out;
SharedReg953_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg953_out;
SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg955_out;
SharedReg1018_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1018_out;
SharedReg909_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg909_out;
SharedReg819_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg819_out;
SharedReg1126_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1126_out;
SharedReg1011_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1011_out;
SharedReg810_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg810_out;
SharedReg540_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg540_out;
SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg326_out;
Delay44No2_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_23_cast <= Delay44No2_out;
Delay45No20_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_24_cast <= Delay45No20_out;
SharedReg958_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg958_out;
SharedReg551_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg551_out;
SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg326_out;
SharedReg811_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg811_out;
   MUX_Subtract18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg539_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg809_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg28_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg472_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg953_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1018_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg909_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg819_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1126_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1011_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg810_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg955_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg540_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay44No2_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay45No20_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg958_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg551_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg326_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg811_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg328_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1014_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg812_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg954_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg18_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg26_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_2_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_2_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Subtract18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Subtract18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Subtract18_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_3_impl_out,
                 X => Delay1No266_out_to_Subtract18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Subtract18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg564_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg564_out;
SharedReg340_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg340_out;
SharedReg553_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg560_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg560_out;
SharedReg557_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg557_out;
SharedReg481_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg481_out;
SharedReg231_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg562_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg1035_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1035_out;
SharedReg664_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg664_out;
SharedReg2_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
SharedReg749_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg749_out;
SharedReg663_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg663_out;
SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg913_out;
SharedReg827_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg827_out;
SharedReg914_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg914_out;
SharedReg828_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg828_out;
SharedReg1025_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1025_out;
SharedReg1136_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1136_out;
SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg556_out;
SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg556_out;
SharedReg128_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg128_out;
SharedReg233_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg233_out;
SharedReg1033_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1033_out;
SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg913_out;
   MUX_Subtract18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg564_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg13_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg10_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg749_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg663_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg827_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg914_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg828_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg553_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1025_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1136_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg556_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg128_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg233_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1033_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg913_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg560_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg557_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg481_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1035_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg664_out_to_MUX_Subtract18_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_3_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_3_impl_0_out,
                 Y => Delay1No266_out);

SharedReg565_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg565_out;
SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg824_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg824_out;
SharedReg553_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg553_out;
SharedReg822_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg822_out;
SharedReg749_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg749_out;
SharedReg340_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg340_out;
SharedReg1027_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1027_out;
SharedReg825_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg825_out;
SharedReg914_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg914_out;
SharedReg18_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
SharedReg478_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg478_out;
SharedReg913_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg913_out;
SharedReg915_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg915_out;
SharedReg1031_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1031_out;
SharedReg900_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg900_out;
SharedReg832_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg832_out;
SharedReg1134_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1134_out;
SharedReg1024_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1024_out;
SharedReg823_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg823_out;
SharedReg554_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg554_out;
SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg338_out;
Delay44No3_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_26_cast <= Delay44No3_out;
Delay45No21_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_27_cast <= Delay45No21_out;
SharedReg918_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg918_out;
   MUX_Subtract18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg565_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg29_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg26_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg478_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg913_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg915_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1031_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg900_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg832_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg824_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1134_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1024_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg823_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg554_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg338_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay44No3_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay45No21_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg918_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg553_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg822_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg749_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg340_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1027_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg825_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg914_out_to_MUX_Subtract18_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_3_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_3_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Subtract18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Subtract18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Subtract18_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_4_impl_out,
                 X => Delay1No268_out_to_Subtract18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Subtract18_4_impl_parent_implementedSystem_port_1_cast);

SharedReg246_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg1046_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1046_out;
SharedReg753_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg753_out;
SharedReg578_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg578_out;
SharedReg352_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg567_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg567_out;
SharedReg574_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg574_out;
SharedReg571_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg571_out;
SharedReg487_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg487_out;
SharedReg244_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg244_out;
SharedReg576_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg576_out;
SharedReg1048_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1048_out;
SharedReg669_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg669_out;
SharedReg2_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg12_out;
SharedReg755_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg755_out;
SharedReg668_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg668_out;
SharedReg903_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg903_out;
SharedReg840_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg840_out;
SharedReg904_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg904_out;
SharedReg841_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg841_out;
SharedReg1038_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1038_out;
SharedReg1144_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1144_out;
SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg570_out;
SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg570_out;
SharedReg138_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg138_out;
   MUX_Subtract18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1046_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg576_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1048_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg669_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg13_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg10_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg12_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg755_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg668_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg903_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg753_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg840_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg904_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg841_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1038_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1144_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg570_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg138_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg578_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg567_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg574_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg571_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg487_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg244_out_to_MUX_Subtract18_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_4_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_4_impl_0_out,
                 Y => Delay1No268_out);

Delay44No4_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_1_cast <= Delay44No4_out;
Delay45No22_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_2_cast <= Delay45No22_out;
SharedReg908_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg579_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg579_out;
SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg350_out;
SharedReg837_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg837_out;
SharedReg567_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg835_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg755_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg755_out;
SharedReg352_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg352_out;
SharedReg1040_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1040_out;
SharedReg838_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg838_out;
SharedReg904_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg904_out;
SharedReg18_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg28_out;
SharedReg484_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg484_out;
SharedReg903_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg903_out;
SharedReg905_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg905_out;
SharedReg1044_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1044_out;
SharedReg453_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg453_out;
SharedReg845_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg845_out;
SharedReg1142_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1142_out;
SharedReg1037_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1037_out;
SharedReg836_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg836_out;
SharedReg568_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg568_out;
SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg350_out;
   MUX_Subtract18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay44No4_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay45No22_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1040_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg838_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg904_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg18_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg29_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg26_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg28_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg484_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg903_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg905_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg908_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1044_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg453_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg845_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1142_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1037_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg836_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg568_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg579_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg350_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg837_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg567_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg755_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg352_out_to_MUX_Subtract18_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_4_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_4_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Subtract18_5_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Subtract18_5_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Subtract18_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_5_impl_out,
                 X => Delay1No270_out_to_Subtract18_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Subtract18_5_impl_parent_implementedSystem_port_1_cast);

SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg584_out;
SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg584_out;
SharedReg148_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg259_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg259_out;
SharedReg1059_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1059_out;
SharedReg932_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg932_out;
SharedReg592_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg592_out;
SharedReg364_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg364_out;
SharedReg581_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg581_out;
SharedReg588_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg588_out;
SharedReg585_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg585_out;
SharedReg493_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg493_out;
SharedReg257_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg257_out;
SharedReg590_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg590_out;
SharedReg1061_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1061_out;
SharedReg674_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg674_out;
SharedReg2_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg12_out;
SharedReg934_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg934_out;
SharedReg673_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg673_out;
SharedReg456_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg456_out;
SharedReg853_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg853_out;
SharedReg457_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg457_out;
SharedReg854_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg854_out;
SharedReg1051_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1051_out;
SharedReg1152_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1152_out;
   MUX_Subtract18_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg584_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg585_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg493_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg257_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg590_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1061_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg674_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg2_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg13_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg10_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg12_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg148_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg934_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg673_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg456_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg853_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg457_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg854_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1051_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1152_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg259_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1059_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg932_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg592_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg364_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg581_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg588_out_to_MUX_Subtract18_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_5_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_5_impl_0_out,
                 Y => Delay1No270_out);

SharedReg849_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg582_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg582_out;
SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg362_out;
Delay44No5_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_4_cast <= Delay44No5_out;
Delay45No23_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_5_cast <= Delay45No23_out;
SharedReg937_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg937_out;
SharedReg593_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg593_out;
SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg850_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg581_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg581_out;
SharedReg848_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg848_out;
SharedReg934_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg934_out;
SharedReg364_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg364_out;
SharedReg1053_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1053_out;
SharedReg851_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg851_out;
SharedReg457_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg457_out;
SharedReg18_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg28_out;
SharedReg490_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg490_out;
SharedReg456_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg456_out;
SharedReg458_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg458_out;
SharedReg1057_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1057_out;
SharedReg440_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg440_out;
SharedReg858_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg858_out;
SharedReg1150_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1150_out;
SharedReg1050_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1050_out;
   MUX_Subtract18_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg582_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg848_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg934_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg364_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1053_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg851_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg457_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg18_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg29_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg26_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg28_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg490_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg456_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg458_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1057_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg440_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg858_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1150_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1050_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => Delay44No5_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay45No23_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg937_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg593_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg581_out_to_MUX_Subtract18_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_5_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_5_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Subtract18_6_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Subtract18_6_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Subtract18_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_6_impl_out,
                 X => Delay1No272_out_to_Subtract18_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Subtract18_6_impl_parent_implementedSystem_port_1_cast);

SharedReg867_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg867_out;
SharedReg1064_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1064_out;
SharedReg1160_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1160_out;
SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg598_out;
SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg598_out;
SharedReg158_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg158_out;
SharedReg272_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg272_out;
SharedReg1072_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1072_out;
SharedReg960_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg960_out;
SharedReg606_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg606_out;
SharedReg376_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg376_out;
SharedReg595_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg595_out;
SharedReg602_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg602_out;
SharedReg599_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg599_out;
SharedReg681_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg681_out;
SharedReg270_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg270_out;
SharedReg604_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg604_out;
SharedReg1074_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1074_out;
SharedReg767_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg767_out;
SharedReg2_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg12_out;
SharedReg962_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg962_out;
SharedReg766_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg766_out;
SharedReg444_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg444_out;
SharedReg866_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg866_out;
SharedReg445_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg445_out;
   MUX_Subtract18_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg867_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1064_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg376_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg595_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg602_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg599_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg681_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg270_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg604_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1074_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg767_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg2_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1160_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg13_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg10_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg12_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg962_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg766_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg444_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg866_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg445_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg598_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg158_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg272_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1072_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg960_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg606_out_to_MUX_Subtract18_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_6_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_6_impl_0_out,
                 Y => Delay1No272_out);

SharedReg871_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg1158_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1158_out;
SharedReg1063_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1063_out;
SharedReg862_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg862_out;
SharedReg596_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg596_out;
SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg374_out;
Delay44No6_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_7_cast <= Delay44No6_out;
Delay45No24_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_8_cast <= Delay45No24_out;
SharedReg925_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg925_out;
SharedReg607_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg607_out;
SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg374_out;
SharedReg863_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg863_out;
SharedReg595_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg595_out;
SharedReg861_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg861_out;
SharedReg962_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg962_out;
SharedReg376_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg376_out;
SharedReg1066_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1066_out;
SharedReg864_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg864_out;
SharedReg445_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg445_out;
SharedReg18_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg28_out;
SharedReg678_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg678_out;
SharedReg444_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg444_out;
SharedReg446_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg446_out;
SharedReg1070_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1070_out;
SharedReg502_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg502_out;
   MUX_Subtract18_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1158_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg863_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg595_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg861_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg962_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg376_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1066_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg864_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg445_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg18_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1063_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg29_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg26_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg28_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg678_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg444_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg446_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1070_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg502_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg862_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg596_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg374_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay44No6_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay45No24_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg925_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg607_out_to_MUX_Subtract18_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_6_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_6_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Subtract18_7_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Subtract18_7_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Subtract18_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_7_impl_out,
                 X => Delay1No274_out_to_Subtract18_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Subtract18_7_impl_parent_implementedSystem_port_1_cast);

SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg966_out;
SharedReg879_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg879_out;
SharedReg967_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg967_out;
SharedReg880_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg880_out;
SharedReg1077_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1077_out;
SharedReg1168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1168_out;
SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg612_out;
SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg612_out;
SharedReg168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg168_out;
SharedReg285_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg285_out;
SharedReg1085_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1085_out;
SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg966_out;
SharedReg620_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg620_out;
SharedReg388_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg388_out;
SharedReg609_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg609_out;
SharedReg616_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg616_out;
SharedReg613_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg613_out;
SharedReg686_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg686_out;
SharedReg283_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg283_out;
SharedReg618_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg618_out;
SharedReg1087_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1087_out;
SharedReg773_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg773_out;
SharedReg2_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg12_out;
SharedReg968_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg968_out;
SharedReg772_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg772_out;
   MUX_Subtract18_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg879_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1085_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg966_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg620_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg388_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg609_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg616_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg613_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg686_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg283_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg618_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg967_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1087_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg773_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg2_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg13_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg10_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg12_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg968_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg772_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg880_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1077_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg612_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg168_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg285_out_to_MUX_Subtract18_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_7_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_7_impl_0_out,
                 Y => Delay1No274_out);

SharedReg639_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg639_out;
SharedReg1083_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1083_out;
SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg637_out;
SharedReg884_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg884_out;
SharedReg1166_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1166_out;
SharedReg1076_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1076_out;
SharedReg875_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg875_out;
SharedReg610_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg610_out;
SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg386_out;
Delay44No7_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_10_cast <= Delay44No7_out;
Delay45No25_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_11_cast <= Delay45No25_out;
SharedReg931_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg931_out;
SharedReg621_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg621_out;
SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg386_out;
SharedReg876_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg876_out;
SharedReg609_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg609_out;
SharedReg874_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg874_out;
SharedReg968_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg968_out;
SharedReg388_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg388_out;
SharedReg1079_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1079_out;
SharedReg877_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg877_out;
SharedReg638_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg638_out;
SharedReg18_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg29_out;
SharedReg26_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg28_out;
SharedReg683_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg683_out;
SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg637_out;
   MUX_Subtract18_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg639_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1083_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay45No25_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg931_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg621_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg876_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg609_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg874_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg968_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg388_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1079_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg877_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg638_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg18_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg29_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg26_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg28_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg683_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg637_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg884_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1166_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1076_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg875_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg610_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg386_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay44No7_out_to_MUX_Subtract18_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_7_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_7_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Subtract18_8_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Subtract18_8_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Subtract18_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_8_impl_out,
                 X => Delay1No276_out_to_Subtract18_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Subtract18_8_impl_parent_implementedSystem_port_1_cast);

SharedReg10_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg780_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg780_out;
SharedReg505_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg505_out;
SharedReg972_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg972_out;
SharedReg892_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg892_out;
SharedReg973_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg973_out;
SharedReg893_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg893_out;
SharedReg1090_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1090_out;
SharedReg1176_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1176_out;
SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg626_out;
SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg626_out;
SharedReg178_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg178_out;
SharedReg298_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg298_out;
SharedReg1098_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1098_out;
SharedReg778_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg778_out;
SharedReg634_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg634_out;
SharedReg400_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg400_out;
SharedReg623_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg623_out;
SharedReg630_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg630_out;
SharedReg627_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg627_out;
SharedReg508_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg508_out;
SharedReg296_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg296_out;
SharedReg632_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg632_out;
SharedReg1100_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1100_out;
SharedReg727_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg727_out;
SharedReg2_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg2_out;
SharedReg13_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg13_out;
   MUX_Subtract18_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg626_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg178_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg298_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1098_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg778_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg634_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg400_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg623_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg630_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg780_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg627_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg508_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg296_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg632_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1100_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg727_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg2_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg13_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg505_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg972_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg892_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg973_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg893_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1090_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1176_out_to_MUX_Subtract18_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_8_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_8_impl_0_out,
                 Y => Delay1No276_out);

SharedReg26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg505_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg505_out;
SharedReg778_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg778_out;
SharedReg974_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg974_out;
SharedReg1096_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1096_out;
SharedReg972_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg972_out;
SharedReg897_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg897_out;
SharedReg1174_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1174_out;
SharedReg1089_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1089_out;
SharedReg888_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg888_out;
SharedReg624_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg624_out;
SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg398_out;
Delay44No8_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_14_cast <= Delay44No8_out;
Delay45No26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_15_cast <= Delay45No26_out;
SharedReg977_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg977_out;
SharedReg635_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg635_out;
SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg398_out;
SharedReg889_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg889_out;
SharedReg623_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg623_out;
SharedReg887_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg887_out;
SharedReg981_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg981_out;
SharedReg400_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg400_out;
SharedReg1092_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1092_out;
SharedReg890_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg890_out;
SharedReg980_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg980_out;
SharedReg18_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg18_out;
SharedReg29_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg29_out;
   MUX_Subtract18_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg888_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg624_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay44No8_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay45No26_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg977_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg635_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg398_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg889_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg623_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg505_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg887_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg981_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg400_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1092_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg890_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg980_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg18_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg29_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg778_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg974_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1096_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg972_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg897_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1174_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1089_out_to_MUX_Subtract18_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract18_8_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_8_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product321_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_0_impl_out,
                 X => Delay1No278_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1275_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1259_out;
SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg1183_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1288_out;
SharedReg1185_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1185_out;
SharedReg305_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg305_out;
SharedReg1187_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1218_out;
SharedReg1236_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1236_out;
SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1110_out;
SharedReg1263_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1263_out;
SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg785_out;
SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg785_out;
SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1112_out;
SharedReg1232_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1232_out;
SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1113_out;
SharedReg1117_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1117_out;
SharedReg1205_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1205_out;
SharedReg1206_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1206_out;
SharedReg41_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg41_out;
SharedReg1207_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1207_out;
   MUX_Product321_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg305_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1187_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1188_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1189_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1218_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1236_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1263_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg785_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1275_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1232_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1113_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1117_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1205_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1206_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg41_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1207_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1281_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1259_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1183_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1288_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1185_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product321_0_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_0_out,
                 Y => Delay1No278_out);

SharedReg1245_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1280_out;
SharedReg1114_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1112_out;
SharedReg1260_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1287_out;
SharedReg185_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg185_out;
SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg987_out;
SharedReg786_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg786_out;
SharedReg1214_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1214_out;
SharedReg516_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg516_out;
SharedReg305_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg305_out;
SharedReg307_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg307_out;
SharedReg37_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg37_out;
SharedReg38_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg38_out;
SharedReg1262_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1262_out;
SharedReg986_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg986_out;
SharedReg1264_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1231_out;
SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg987_out;
SharedReg1233_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1233_out;
SharedReg1237_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1237_out;
SharedReg199_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg199_out;
SharedReg40_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg40_out;
SharedReg1234_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1234_out;
SharedReg39_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg39_out;
   MUX_Product321_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1245_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1280_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1214_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg516_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg305_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg307_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg37_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg38_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1262_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg986_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1264_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1265_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1231_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1233_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1237_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg199_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg40_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1234_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg39_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1112_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1260_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1287_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg185_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg987_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg786_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product321_0_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product321_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_1_impl_out,
                 X => Delay1No280_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1206_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1206_out;
SharedReg48_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg1207_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1207_out;
SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1118_out;
SharedReg1121_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1121_out;
SharedReg1275_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1275_out;
SharedReg1281_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1281_out;
SharedReg1259_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1259_out;
SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1120_out;
SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg1183_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1183_out;
SharedReg1288_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1288_out;
SharedReg1185_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1185_out;
SharedReg317_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg317_out;
SharedReg1187_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1187_out;
SharedReg1188_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1188_out;
SharedReg1189_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1189_out;
SharedReg1218_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1218_out;
SharedReg1236_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1236_out;
SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1118_out;
SharedReg1263_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1263_out;
SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg798_out;
SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg798_out;
SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1120_out;
SharedReg1202_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1202_out;
SharedReg1203_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1203_out;
SharedReg1204_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1204_out;
SharedReg212_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg212_out;
   MUX_Product321_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1206_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1183_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1288_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1185_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg317_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1187_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1188_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1189_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1218_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1236_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1207_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1263_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg798_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1202_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1203_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1204_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg212_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1121_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1275_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1281_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1259_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1120_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product321_1_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_0_out,
                 Y => Delay1No280_out);

SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg1234_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1234_out;
SharedReg46_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg1245_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1245_out;
SharedReg1280_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1280_out;
SharedReg1122_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1122_out;
SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1120_out;
SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1260_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1260_out;
SharedReg1287_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1287_out;
SharedReg198_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg198_out;
SharedReg1000_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1000_out;
SharedReg799_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg799_out;
SharedReg1214_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1214_out;
SharedReg530_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg530_out;
SharedReg317_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg317_out;
SharedReg319_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg319_out;
SharedReg44_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg44_out;
SharedReg45_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg45_out;
SharedReg1262_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1262_out;
SharedReg999_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg999_out;
SharedReg1264_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1265_out;
SharedReg1231_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1231_out;
SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg47_out;
SharedReg115_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg115_out;
SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg47_out;
SharedReg1232_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1232_out;
   MUX_Product321_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1234_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg198_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1000_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg799_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1214_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg530_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg317_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg319_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg44_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg45_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1262_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg46_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg999_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1264_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1265_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1231_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg115_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg47_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1232_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg1245_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1280_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1122_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1260_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1287_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Product321_1_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Subtract22_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_0_impl_out,
                 X => Delay1No282_out_to_Subtract22_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Subtract22_0_impl_parent_implementedSystem_port_1_cast);

SharedReg648_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg648_out;
SharedReg3_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg733_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg733_out;
SharedReg736_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg736_out;
SharedReg515_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg515_out;
SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg189_out;
SharedReg516_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg516_out;
SharedReg307_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg307_out;
SharedReg186_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg186_out;
SharedReg304_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg304_out;
SharedReg34_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg34_out;
SharedReg185_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg185_out;
SharedReg512_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg512_out;
SharedReg1102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1102_out;
SharedReg194_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg194_out;
SharedReg517_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg517_out;
SharedReg102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg102_out;
SharedReg1116_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1116_out;
SharedReg302_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg302_out;
SharedReg306_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg306_out;
SharedReg101_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg101_out;
SharedReg785_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg785_out;
SharedReg790_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg790_out;
SharedReg192_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg192_out;
SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg195_out;
   MUX_Subtract22_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg648_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg307_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg186_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg304_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg34_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg185_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg512_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg194_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg517_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg102_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg15_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1116_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg302_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg306_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg101_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg785_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg790_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg192_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg195_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg11_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg733_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg736_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg515_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg189_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg516_out_to_MUX_Subtract22_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_0_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_0_impl_0_out,
                 Y => Delay1No282_out);

SharedReg939_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg939_out;
SharedReg19_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1103_out;
SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1103_out;
SharedReg519_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg519_out;
SharedReg308_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg308_out;
SharedReg521_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg309_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg309_out;
SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg302_out;
SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg302_out;
SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg302_out;
SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg302_out;
SharedReg986_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg986_out;
SharedReg1104_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1104_out;
SharedReg197_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg197_out;
SharedReg787_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg787_out;
SharedReg196_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg196_out;
SharedReg794_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg794_out;
SharedReg304_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg304_out;
SharedReg95_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg95_out;
SharedReg185_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg185_out;
SharedReg1113_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1113_out;
SharedReg512_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg512_out;
SharedReg35_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg35_out;
SharedReg305_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg305_out;
   MUX_Subtract22_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg939_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg309_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg302_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg986_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1104_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg197_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg787_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg196_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg31_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg794_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg304_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg95_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg185_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1113_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg512_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg35_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg305_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg27_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1103_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg519_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg308_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Subtract22_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_0_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_0_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Subtract22_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_1_impl_out,
                 X => Delay1No284_out_to_Subtract22_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Subtract22_1_impl_parent_implementedSystem_port_1_cast);

SharedReg803_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg205_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg208_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg208_out;
SharedReg466_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg466_out;
SharedReg3_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg14_out;
SharedReg738_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg738_out;
SharedReg741_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg741_out;
SharedReg529_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg529_out;
SharedReg202_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg202_out;
SharedReg530_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg530_out;
SharedReg319_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg319_out;
SharedReg199_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg199_out;
SharedReg316_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg316_out;
SharedReg41_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg41_out;
SharedReg198_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg198_out;
SharedReg526_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg526_out;
SharedReg1106_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1106_out;
SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg207_out;
SharedReg531_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg531_out;
SharedReg112_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg112_out;
SharedReg1124_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1124_out;
SharedReg314_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg314_out;
SharedReg318_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg318_out;
SharedReg111_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg111_out;
SharedReg798_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg798_out;
   MUX_Subtract22_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg529_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg530_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg319_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg199_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg316_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg41_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg198_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg526_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1106_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg208_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg207_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg531_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg112_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1124_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg314_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg318_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg111_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg798_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg466_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg14_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg738_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg741_out_to_MUX_Subtract22_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_1_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_1_impl_0_out,
                 Y => Delay1No284_out);

SharedReg526_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg526_out;
SharedReg42_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg317_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg737_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg737_out;
SharedReg19_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1107_out;
SharedReg533_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg533_out;
SharedReg320_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg320_out;
SharedReg535_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg535_out;
SharedReg321_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg321_out;
SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg314_out;
SharedReg999_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg999_out;
SharedReg1108_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1108_out;
SharedReg210_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg210_out;
SharedReg800_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg800_out;
SharedReg209_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg209_out;
SharedReg807_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg807_out;
SharedReg316_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg316_out;
SharedReg105_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg105_out;
SharedReg198_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg198_out;
SharedReg1121_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1121_out;
   MUX_Subtract22_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg526_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg533_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg320_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg535_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg321_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg314_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg999_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1108_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg317_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg210_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg800_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg209_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg807_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg316_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg105_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg198_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1121_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg737_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1107_out_to_MUX_Subtract22_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_1_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_1_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Subtract22_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_2_impl_out,
                 X => Delay1No286_out_to_Subtract22_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Subtract22_2_impl_parent_implementedSystem_port_1_cast);

SharedReg330_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg330_out;
SharedReg121_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg811_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg811_out;
SharedReg816_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg218_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg221_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg221_out;
SharedReg472_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg472_out;
SharedReg3_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg14_out;
SharedReg743_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg743_out;
SharedReg746_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg746_out;
SharedReg543_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg543_out;
SharedReg215_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg215_out;
SharedReg544_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg544_out;
SharedReg331_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg331_out;
SharedReg212_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg212_out;
SharedReg328_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg328_out;
SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg48_out;
SharedReg211_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg211_out;
SharedReg540_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg540_out;
SharedReg909_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg909_out;
SharedReg220_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg220_out;
SharedReg545_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg545_out;
SharedReg122_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg122_out;
SharedReg1132_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1132_out;
SharedReg326_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg326_out;
   MUX_Subtract22_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg330_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg14_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg743_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg746_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg543_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg215_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg544_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg331_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg212_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg328_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg48_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg811_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg211_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg540_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg909_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg220_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg545_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg122_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1132_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg326_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg816_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg221_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg472_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg15_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Subtract22_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_2_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_2_impl_0_out,
                 Y => Delay1No286_out);

SharedReg115_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg211_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg1129_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1129_out;
SharedReg540_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg540_out;
SharedReg49_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg49_out;
SharedReg329_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg329_out;
SharedReg742_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg742_out;
SharedReg19_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg30_out;
SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg910_out;
SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg910_out;
SharedReg547_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg547_out;
SharedReg332_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg332_out;
SharedReg549_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg549_out;
SharedReg333_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg333_out;
SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg326_out;
SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg326_out;
SharedReg1012_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1012_out;
SharedReg911_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg911_out;
SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg223_out;
SharedReg813_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg813_out;
SharedReg222_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg222_out;
SharedReg820_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg820_out;
SharedReg328_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg328_out;
   MUX_Subtract22_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg30_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg910_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg547_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg332_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg549_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg333_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1129_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg326_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1012_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg911_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg223_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg813_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg222_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg820_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg328_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg540_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg49_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg329_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg742_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Subtract22_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_2_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_2_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Subtract22_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_3_impl_out,
                 X => Delay1No288_out_to_Subtract22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Subtract22_3_impl_parent_implementedSystem_port_1_cast);

SharedReg132_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg1140_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1140_out;
SharedReg338_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg342_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg342_out;
SharedReg131_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg131_out;
SharedReg824_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg824_out;
SharedReg829_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg231_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg231_out;
SharedReg234_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg234_out;
SharedReg478_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg478_out;
SharedReg3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg14_out;
SharedReg748_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg748_out;
SharedReg751_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg751_out;
SharedReg557_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg557_out;
SharedReg228_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg228_out;
SharedReg558_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg558_out;
SharedReg343_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg343_out;
SharedReg225_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg225_out;
SharedReg340_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg340_out;
SharedReg55_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg55_out;
SharedReg224_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg224_out;
SharedReg554_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg554_out;
SharedReg900_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg900_out;
SharedReg233_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg233_out;
SharedReg559_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg559_out;
   MUX_Subtract22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1140_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg15_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg11_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg14_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg748_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg751_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg557_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg228_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg558_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg343_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg338_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg225_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg340_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg55_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg224_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg554_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg900_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg233_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg559_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg342_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg131_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg824_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg231_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg234_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg478_out_to_MUX_Subtract22_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_3_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_3_impl_0_out,
                 Y => Delay1No288_out);

SharedReg235_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg833_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg833_out;
SharedReg340_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg340_out;
SharedReg125_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg125_out;
SharedReg224_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg1137_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1137_out;
SharedReg554_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg554_out;
SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg56_out;
SharedReg341_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg341_out;
SharedReg747_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg747_out;
SharedReg19_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg901_out;
SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg901_out;
SharedReg561_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg561_out;
SharedReg344_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg344_out;
SharedReg563_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg563_out;
SharedReg345_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg345_out;
SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg338_out;
SharedReg1025_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1025_out;
SharedReg902_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg902_out;
SharedReg236_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg236_out;
SharedReg826_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg826_out;
   MUX_Subtract22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg833_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg27_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg901_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg561_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg344_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg563_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg345_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg340_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg338_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1025_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg902_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg236_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg826_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg125_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1137_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg554_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg56_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg341_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg747_out_to_MUX_Subtract22_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_3_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_3_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Subtract22_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_4_impl_out,
                 X => Delay1No290_out_to_Subtract22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Subtract22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg246_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg246_out;
SharedReg573_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg573_out;
SharedReg142_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg142_out;
SharedReg1148_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1148_out;
SharedReg350_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg350_out;
SharedReg354_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg354_out;
SharedReg141_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg141_out;
SharedReg837_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg842_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg842_out;
SharedReg244_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg244_out;
SharedReg247_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg247_out;
SharedReg484_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg484_out;
SharedReg3_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg14_out;
SharedReg754_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg754_out;
SharedReg757_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg757_out;
SharedReg571_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg571_out;
SharedReg241_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg241_out;
SharedReg572_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg572_out;
SharedReg355_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg355_out;
SharedReg238_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg238_out;
SharedReg352_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg352_out;
SharedReg62_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg62_out;
SharedReg237_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg237_out;
SharedReg568_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg568_out;
   MUX_Subtract22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg246_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg244_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg247_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg484_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg3_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg15_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg11_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg14_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg754_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg757_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg571_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg573_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg241_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg572_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg355_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg238_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg352_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg62_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg237_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg568_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg142_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1148_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg354_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg141_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg842_out_to_MUX_Subtract22_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_4_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_4_impl_0_out,
                 Y => Delay1No290_out);

SharedReg455_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg455_out;
SharedReg249_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg839_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg839_out;
SharedReg248_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg248_out;
SharedReg846_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg846_out;
SharedReg352_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg352_out;
SharedReg135_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg135_out;
SharedReg237_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg237_out;
SharedReg1145_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1145_out;
SharedReg568_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg63_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg63_out;
SharedReg353_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg353_out;
SharedReg753_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg753_out;
SharedReg19_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg30_out;
SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg454_out;
SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg454_out;
SharedReg575_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg575_out;
SharedReg356_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg356_out;
SharedReg577_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg577_out;
SharedReg357_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg357_out;
SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg350_out;
SharedReg1038_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1038_out;
   MUX_Subtract22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg455_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg63_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg353_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg753_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg19_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg31_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg27_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg30_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg454_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg575_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg839_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg356_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg577_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg357_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg350_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1038_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg248_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg846_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg352_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg135_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg237_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1145_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Subtract22_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_4_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_4_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Subtract22_5_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Subtract22_5_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Subtract22_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_5_impl_out,
                 X => Delay1No292_out_to_Subtract22_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Subtract22_5_impl_parent_implementedSystem_port_1_cast);

SharedReg69_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg250_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg250_out;
SharedReg582_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg582_out;
SharedReg932_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg932_out;
SharedReg259_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg259_out;
SharedReg587_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg587_out;
SharedReg152_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg152_out;
SharedReg1156_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1156_out;
SharedReg362_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg362_out;
SharedReg366_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg366_out;
SharedReg151_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg850_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg850_out;
SharedReg855_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg855_out;
SharedReg257_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg257_out;
SharedReg260_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg260_out;
SharedReg490_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg490_out;
SharedReg3_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg14_out;
SharedReg933_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg933_out;
SharedReg936_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg936_out;
SharedReg585_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg585_out;
SharedReg254_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg254_out;
SharedReg586_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg586_out;
SharedReg367_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg367_out;
SharedReg251_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg251_out;
SharedReg364_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg364_out;
   MUX_Subtract22_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg250_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg850_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg855_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg257_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg260_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg490_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg3_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg15_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg11_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg14_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg582_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg933_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg936_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg585_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg254_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg586_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg367_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg251_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg364_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg932_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg587_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg152_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1156_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg362_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg366_out_to_MUX_Subtract22_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_5_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_5_impl_0_out,
                 Y => Delay1No292_out);

SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg362_out;
SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg362_out;
SharedReg1051_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1051_out;
SharedReg458_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg458_out;
SharedReg262_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg852_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg852_out;
SharedReg261_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg859_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg859_out;
SharedReg364_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg364_out;
SharedReg145_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg145_out;
SharedReg250_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg250_out;
SharedReg1153_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1153_out;
SharedReg582_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg582_out;
SharedReg70_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg70_out;
SharedReg365_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg365_out;
SharedReg932_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg932_out;
SharedReg19_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg30_out;
SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg441_out;
SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg441_out;
SharedReg589_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg589_out;
SharedReg368_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg368_out;
SharedReg591_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg591_out;
SharedReg369_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg369_out;
SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg362_out;
SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg362_out;
   MUX_Subtract22_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1153_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg582_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg70_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg365_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg932_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg19_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg31_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg27_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg30_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1051_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg441_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg589_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg368_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg591_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg369_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg362_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg458_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg852_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg859_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg364_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg145_out_to_MUX_Subtract22_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_5_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_5_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Subtract22_6_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Subtract22_6_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Subtract22_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_6_impl_out,
                 X => Delay1No294_out_to_Subtract22_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Subtract22_6_impl_parent_implementedSystem_port_1_cast);

SharedReg379_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg264_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg376_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg376_out;
SharedReg76_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg76_out;
SharedReg263_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg263_out;
SharedReg596_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg596_out;
SharedReg960_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg960_out;
SharedReg272_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg272_out;
SharedReg601_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg601_out;
SharedReg162_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg162_out;
SharedReg1164_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1164_out;
SharedReg374_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg374_out;
SharedReg378_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg378_out;
SharedReg161_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg161_out;
SharedReg863_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg863_out;
SharedReg868_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg868_out;
SharedReg270_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg270_out;
SharedReg273_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg273_out;
SharedReg678_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg678_out;
SharedReg3_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg14_out;
SharedReg961_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg961_out;
SharedReg964_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg964_out;
SharedReg599_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg599_out;
SharedReg267_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg267_out;
SharedReg600_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg600_out;
   MUX_Subtract22_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1164_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg374_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg378_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg161_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg863_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg868_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg270_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg273_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg678_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg3_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg376_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg15_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg11_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg14_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg961_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg964_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg599_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg267_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg600_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg76_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg263_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg596_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg960_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg272_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg601_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg162_out_to_MUX_Subtract22_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_6_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_6_impl_0_out,
                 Y => Delay1No294_out);

SharedReg381_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg381_out;
SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg374_out;
SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg374_out;
SharedReg1064_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1064_out;
SharedReg446_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg446_out;
SharedReg275_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg275_out;
SharedReg865_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg865_out;
SharedReg274_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg274_out;
SharedReg872_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg872_out;
SharedReg376_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg376_out;
SharedReg155_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg155_out;
SharedReg263_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg263_out;
SharedReg1161_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1161_out;
SharedReg596_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg596_out;
SharedReg77_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg77_out;
SharedReg377_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg377_out;
SharedReg960_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg960_out;
SharedReg19_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg30_out;
SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg503_out;
SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg503_out;
SharedReg603_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg603_out;
SharedReg380_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg380_out;
SharedReg605_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg605_out;
   MUX_Subtract22_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg381_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg872_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg376_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg155_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg263_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1161_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg596_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg77_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg377_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg960_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg19_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg31_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg27_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg30_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg503_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg603_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg380_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg605_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg374_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1064_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg446_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg275_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg865_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg274_out_to_MUX_Subtract22_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_6_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_6_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Subtract22_7_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Subtract22_7_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Subtract22_7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_7_impl_out,
                 X => Delay1No296_out_to_Subtract22_7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Subtract22_7_impl_parent_implementedSystem_port_1_cast);

SharedReg613_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg613_out;
SharedReg280_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
SharedReg614_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg614_out;
SharedReg391_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg391_out;
SharedReg277_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_5_cast <= SharedReg277_out;
SharedReg388_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_6_cast <= SharedReg388_out;
SharedReg83_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_7_cast <= SharedReg83_out;
SharedReg276_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_8_cast <= SharedReg276_out;
SharedReg610_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_9_cast <= SharedReg610_out;
SharedReg966_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_10_cast <= SharedReg966_out;
SharedReg285_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_11_cast <= SharedReg285_out;
SharedReg615_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_12_cast <= SharedReg615_out;
SharedReg172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_13_cast <= SharedReg172_out;
SharedReg1172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1172_out;
SharedReg386_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_15_cast <= SharedReg386_out;
SharedReg390_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_16_cast <= SharedReg390_out;
SharedReg171_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_17_cast <= SharedReg171_out;
SharedReg876_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_18_cast <= SharedReg876_out;
SharedReg881_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_19_cast <= SharedReg881_out;
SharedReg283_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_20_cast <= SharedReg283_out;
SharedReg286_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_21_cast <= SharedReg286_out;
SharedReg683_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_22_cast <= SharedReg683_out;
SharedReg3_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_23_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_24_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_25_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_26_cast <= SharedReg14_out;
SharedReg967_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_27_cast <= SharedReg967_out;
SharedReg970_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_28_cast <= SharedReg970_out;
   MUX_Subtract22_7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg613_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg285_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg615_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1172_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg386_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg390_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg171_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg876_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg881_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg283_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg614_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg286_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg683_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg3_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg15_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg11_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg14_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg967_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg970_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg391_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg277_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg388_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg83_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg276_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg610_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg966_out_to_MUX_Subtract22_7_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_7_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_7_impl_0_out,
                 Y => Delay1No296_out);

SharedReg617_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg617_out;
SharedReg392_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg619_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg619_out;
SharedReg393_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg393_out;
SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_5_cast <= SharedReg386_out;
SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_6_cast <= SharedReg386_out;
SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_8_cast <= SharedReg386_out;
SharedReg1077_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1077_out;
SharedReg639_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_10_cast <= SharedReg639_out;
SharedReg288_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_11_cast <= SharedReg288_out;
SharedReg878_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_12_cast <= SharedReg878_out;
SharedReg287_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_13_cast <= SharedReg287_out;
SharedReg885_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_14_cast <= SharedReg885_out;
SharedReg388_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_15_cast <= SharedReg388_out;
SharedReg165_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_16_cast <= SharedReg165_out;
SharedReg276_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_17_cast <= SharedReg276_out;
SharedReg1169_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1169_out;
SharedReg610_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_19_cast <= SharedReg610_out;
SharedReg84_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_20_cast <= SharedReg84_out;
SharedReg389_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_21_cast <= SharedReg389_out;
SharedReg966_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_22_cast <= SharedReg966_out;
SharedReg19_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_23_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_24_cast <= SharedReg31_out;
SharedReg27_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_25_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_26_cast <= SharedReg30_out;
SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_27_cast <= SharedReg451_out;
SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_28_cast <= SharedReg451_out;
   MUX_Subtract22_7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg617_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg288_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg878_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg287_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg885_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg388_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg165_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg276_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1169_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg610_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg84_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg619_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg389_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg966_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg19_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg31_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg27_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg30_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg451_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg393_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg386_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1077_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg639_out_to_MUX_Subtract22_7_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_7_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_7_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Subtract22_8_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Subtract22_8_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Subtract22_8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_8_impl_out,
                 X => Delay1No298_out_to_Subtract22_8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Subtract22_8_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg14_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg779_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg779_out;
SharedReg976_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg976_out;
SharedReg627_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg293_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_6_cast <= SharedReg293_out;
SharedReg628_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_7_cast <= SharedReg628_out;
SharedReg403_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_8_cast <= SharedReg403_out;
SharedReg290_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_9_cast <= SharedReg290_out;
SharedReg400_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_10_cast <= SharedReg400_out;
SharedReg90_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_11_cast <= SharedReg90_out;
SharedReg289_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_12_cast <= SharedReg289_out;
SharedReg624_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_13_cast <= SharedReg624_out;
SharedReg979_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_14_cast <= SharedReg979_out;
SharedReg298_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_15_cast <= SharedReg298_out;
SharedReg629_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_16_cast <= SharedReg629_out;
SharedReg182_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_17_cast <= SharedReg182_out;
SharedReg1180_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1180_out;
SharedReg398_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_19_cast <= SharedReg398_out;
SharedReg402_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_20_cast <= SharedReg402_out;
SharedReg181_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_21_cast <= SharedReg181_out;
SharedReg889_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_22_cast <= SharedReg889_out;
SharedReg894_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_23_cast <= SharedReg894_out;
SharedReg296_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_24_cast <= SharedReg296_out;
SharedReg299_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_25_cast <= SharedReg299_out;
SharedReg726_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_26_cast <= SharedReg726_out;
SharedReg3_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_27_cast <= SharedReg3_out;
SharedReg15_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_28_cast <= SharedReg15_out;
   MUX_Subtract22_8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg90_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg289_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg624_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg979_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg298_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg629_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg182_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1180_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg398_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg402_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg779_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg181_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg889_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg894_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg296_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg299_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg726_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg3_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg15_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg976_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg293_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg628_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg403_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg290_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg400_out_to_MUX_Subtract22_8_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_8_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_8_impl_0_out,
                 Y => Delay1No298_out);

SharedReg27_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg30_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg980_out;
SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg980_out;
SharedReg631_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_5_cast <= SharedReg631_out;
SharedReg404_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg633_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_7_cast <= SharedReg633_out;
SharedReg405_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_8_cast <= SharedReg405_out;
SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_9_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_10_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_11_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_12_cast <= SharedReg398_out;
SharedReg1090_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1090_out;
SharedReg981_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_14_cast <= SharedReg981_out;
SharedReg301_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_15_cast <= SharedReg301_out;
SharedReg891_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_16_cast <= SharedReg891_out;
SharedReg300_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_17_cast <= SharedReg300_out;
SharedReg898_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_18_cast <= SharedReg898_out;
SharedReg400_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_19_cast <= SharedReg400_out;
SharedReg175_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_20_cast <= SharedReg175_out;
SharedReg289_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_21_cast <= SharedReg289_out;
SharedReg1177_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1177_out;
SharedReg624_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_23_cast <= SharedReg624_out;
SharedReg91_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_24_cast <= SharedReg91_out;
SharedReg401_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_25_cast <= SharedReg401_out;
SharedReg979_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_26_cast <= SharedReg979_out;
SharedReg19_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_27_cast <= SharedReg19_out;
SharedReg31_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_28_cast <= SharedReg31_out;
   MUX_Subtract22_8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_28_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1090_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg981_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg301_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg891_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg300_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg898_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg400_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg175_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg289_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1177_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg624_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg91_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg401_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg979_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg19_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg31_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_28_cast,
                 iS_3 => SharedReg980_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg631_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg633_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg405_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg398_out_to_MUX_Subtract22_8_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount281_out,
                 oMux => MUX_Subtract22_8_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_8_impl_1_out,
                 Y => Delay1No299_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay4No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => Delay4No233_out);

   Delay4No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => Delay4No241_out);

   Delay8No27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => Delay8No27_out);

   Delay8No28_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => Delay8No28_out);

   Delay8No29_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => Delay8No29_out);

   Delay8No30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => Delay8No30_out);

   Delay8No31_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => Delay8No31_out);

   Delay8No32_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => Delay8No32_out);

   Delay8No33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => Delay8No33_out);

   Delay8No34_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => Delay8No34_out);

   Delay8No35_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => Delay8No35_out);

   Delay8No36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => Delay8No36_out);

   Delay8No37_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => Delay8No37_out);

   Delay8No38_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => Delay8No38_out);

   Delay8No39_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => Delay8No39_out);

   Delay8No42_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => Delay8No42_out);

   Delay8No43_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => Delay8No43_out);

   Delay8No44_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => Delay8No44_out);

   Delay6No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => Delay6No90_out);

   Delay6No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => Delay6No91_out);

   Delay6No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => Delay6No92_out);

   Delay6No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => Delay6No93_out);

   Delay6No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => Delay6No94_out);

   Delay6No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => Delay6No95_out);

   Delay6No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => Delay6No105_out);

   Delay6No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => Delay6No108_out);

   Delay6No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => Delay6No109_out);

   Delay6No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => Delay6No110_out);

   Delay6No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => Delay6No111_out);

   Delay6No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => Delay6No112_out);

   Delay6No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => Delay6No113_out);

   Delay6No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => Delay6No125_out);

   Delay9No18_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => Delay9No18_out);

   Delay9No19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => Delay9No19_out);

   Delay9No20_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => Delay9No20_out);

   Delay9No31_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => Delay9No31_out);

   Delay9No32_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => Delay9No32_out);

   Delay9No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => Delay9No33_out);

   Delay9No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => Delay9No34_out);

   Delay10No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => Delay10No18_out);

   Delay10No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => Delay10No19_out);

   Delay10No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => Delay10No20_out);

   Delay10No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => Delay10No21_out);

   Delay10No22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => Delay10No22_out);

   Delay10No23_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => Delay10No23_out);

   Delay10No24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => Delay10No24_out);

   Delay10No25_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => Delay10No25_out);

   Delay10No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => Delay10No26_out);

   Delay9No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1105_out,
                 Y => Delay9No36_out);

   Delay9No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1109_out,
                 Y => Delay9No37_out);

   Delay9No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => Delay9No38_out);

   Delay44No_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => Delay44No_out);

   Delay44No1_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => Delay44No1_out);

   Delay44No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => Delay44No2_out);

   Delay44No3_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => Delay44No3_out);

   Delay44No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => Delay44No4_out);

   Delay44No5_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => Delay44No5_out);

   Delay44No6_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => Delay44No6_out);

   Delay44No7_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => Delay44No7_out);

   Delay44No8_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => Delay44No8_out);

   Delay45No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => Delay45No18_out);

   Delay45No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => Delay45No19_out);

   Delay45No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => Delay45No20_out);

   Delay45No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => Delay45No21_out);

   Delay45No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => Delay45No22_out);

   Delay45No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => Delay45No23_out);

   Delay45No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => Delay45No24_out);

   Delay45No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => Delay45No25_out);

   Delay45No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => Delay45No26_out);

   Delay27No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => Delay27No_out);

   Delay27No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay27No1_out);

   Delay27No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => Delay27No2_out);

   Delay27No3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => Delay27No3_out);

   Delay27No4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => Delay27No4_out);

   Delay27No5_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => Delay27No5_out);

   Delay27No6_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => Delay27No6_out);

   Delay27No7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => Delay27No7_out);

   Delay27No8_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay27No8_out);

   Delay8No111_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => Delay8No111_out);

   Delay8No112_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => Delay8No112_out);

   Delay8No113_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => Delay8No113_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_5_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Product316_8_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product316_8_impl_0_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product316_8_impl_0_LUT_out);

   MUX_Product316_8_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product316_8_impl_1_LUT_wIn_5_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount281_out,
                 Output => MUX_Product316_8_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_5_impl_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_6_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_7_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_8_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_5_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_6_impl_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_7_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_8_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_0_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_1_impl_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_2_impl_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_3_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_4_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_5_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_6_impl_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_7_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_8_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_2_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_3_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_4_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_5_impl_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_6_impl_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_7_impl_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_8_impl_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_5_impl_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_6_impl_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_7_impl_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_8_impl_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_5_impl_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_6_impl_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_4_impl_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_5_impl_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_6_impl_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_7_impl_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_8_impl_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_5_impl_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_6_impl_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_7_impl_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_8_impl_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_8_impl_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_7_impl_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_5_impl_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_6_impl_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_7_impl_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_8_impl_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_0_impl_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_1_impl_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_2_impl_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_3_impl_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_4_impl_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_8_impl_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_0_impl_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_1_impl_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_2_impl_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_3_impl_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_4_impl_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_5_impl_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_6_impl_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_7_impl_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_8_impl_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_0_impl_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_2_impl_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_3_impl_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_4_impl_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_5_impl_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg857_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_6_impl_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_7_impl_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_8_impl_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product34_4_impl_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product34_5_impl_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_3_impl_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_4_impl_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg918_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_6_impl_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_7_impl_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_5_impl_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg934_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_0_impl_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_1_impl_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_2_impl_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_6_impl_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_7_impl_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg967_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_8_impl_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product316_8_impl_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg983_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_0_impl_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg985_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_1_impl_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1000_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1003_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1006_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_2_impl_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);

   SharedReg1015_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => SharedReg1015_out);

   SharedReg1016_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1015_out,
                 Y => SharedReg1016_out);

   SharedReg1017_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1016_out,
                 Y => SharedReg1017_out);

   SharedReg1018_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1017_out,
                 Y => SharedReg1018_out);

   SharedReg1019_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1018_out,
                 Y => SharedReg1019_out);

   SharedReg1020_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1019_out,
                 Y => SharedReg1020_out);

   SharedReg1021_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1020_out,
                 Y => SharedReg1021_out);

   SharedReg1022_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1021_out,
                 Y => SharedReg1022_out);

   SharedReg1023_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1022_out,
                 Y => SharedReg1023_out);

   SharedReg1024_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_3_impl_out,
                 Y => SharedReg1024_out);

   SharedReg1025_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1024_out,
                 Y => SharedReg1025_out);

   SharedReg1026_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1025_out,
                 Y => SharedReg1026_out);

   SharedReg1027_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1026_out,
                 Y => SharedReg1027_out);

   SharedReg1028_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1027_out,
                 Y => SharedReg1028_out);

   SharedReg1029_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1028_out,
                 Y => SharedReg1029_out);

   SharedReg1030_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1029_out,
                 Y => SharedReg1030_out);

   SharedReg1031_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1030_out,
                 Y => SharedReg1031_out);

   SharedReg1032_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1031_out,
                 Y => SharedReg1032_out);

   SharedReg1033_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1032_out,
                 Y => SharedReg1033_out);

   SharedReg1034_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1033_out,
                 Y => SharedReg1034_out);

   SharedReg1035_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1034_out,
                 Y => SharedReg1035_out);

   SharedReg1036_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1035_out,
                 Y => SharedReg1036_out);

   SharedReg1037_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_4_impl_out,
                 Y => SharedReg1037_out);

   SharedReg1038_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1037_out,
                 Y => SharedReg1038_out);

   SharedReg1039_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1038_out,
                 Y => SharedReg1039_out);

   SharedReg1040_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1039_out,
                 Y => SharedReg1040_out);

   SharedReg1041_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1040_out,
                 Y => SharedReg1041_out);

   SharedReg1042_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1041_out,
                 Y => SharedReg1042_out);

   SharedReg1043_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1042_out,
                 Y => SharedReg1043_out);

   SharedReg1044_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1043_out,
                 Y => SharedReg1044_out);

   SharedReg1045_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1044_out,
                 Y => SharedReg1045_out);

   SharedReg1046_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1045_out,
                 Y => SharedReg1046_out);

   SharedReg1047_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1046_out,
                 Y => SharedReg1047_out);

   SharedReg1048_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1047_out,
                 Y => SharedReg1048_out);

   SharedReg1049_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1048_out,
                 Y => SharedReg1049_out);

   SharedReg1050_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_5_impl_out,
                 Y => SharedReg1050_out);

   SharedReg1051_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1050_out,
                 Y => SharedReg1051_out);

   SharedReg1052_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1051_out,
                 Y => SharedReg1052_out);

   SharedReg1053_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1052_out,
                 Y => SharedReg1053_out);

   SharedReg1054_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1053_out,
                 Y => SharedReg1054_out);

   SharedReg1055_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1054_out,
                 Y => SharedReg1055_out);

   SharedReg1056_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1055_out,
                 Y => SharedReg1056_out);

   SharedReg1057_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1056_out,
                 Y => SharedReg1057_out);

   SharedReg1058_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1057_out,
                 Y => SharedReg1058_out);

   SharedReg1059_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1058_out,
                 Y => SharedReg1059_out);

   SharedReg1060_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1059_out,
                 Y => SharedReg1060_out);

   SharedReg1061_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1060_out,
                 Y => SharedReg1061_out);

   SharedReg1062_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1061_out,
                 Y => SharedReg1062_out);

   SharedReg1063_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_6_impl_out,
                 Y => SharedReg1063_out);

   SharedReg1064_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1063_out,
                 Y => SharedReg1064_out);

   SharedReg1065_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1064_out,
                 Y => SharedReg1065_out);

   SharedReg1066_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1065_out,
                 Y => SharedReg1066_out);

   SharedReg1067_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1066_out,
                 Y => SharedReg1067_out);

   SharedReg1068_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1067_out,
                 Y => SharedReg1068_out);

   SharedReg1069_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1068_out,
                 Y => SharedReg1069_out);

   SharedReg1070_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1069_out,
                 Y => SharedReg1070_out);

   SharedReg1071_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1070_out,
                 Y => SharedReg1071_out);

   SharedReg1072_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1071_out,
                 Y => SharedReg1072_out);

   SharedReg1073_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1072_out,
                 Y => SharedReg1073_out);

   SharedReg1074_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1073_out,
                 Y => SharedReg1074_out);

   SharedReg1075_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1074_out,
                 Y => SharedReg1075_out);

   SharedReg1076_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_7_impl_out,
                 Y => SharedReg1076_out);

   SharedReg1077_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1076_out,
                 Y => SharedReg1077_out);

   SharedReg1078_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1077_out,
                 Y => SharedReg1078_out);

   SharedReg1079_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1078_out,
                 Y => SharedReg1079_out);

   SharedReg1080_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1079_out,
                 Y => SharedReg1080_out);

   SharedReg1081_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1080_out,
                 Y => SharedReg1081_out);

   SharedReg1082_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1081_out,
                 Y => SharedReg1082_out);

   SharedReg1083_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1082_out,
                 Y => SharedReg1083_out);

   SharedReg1084_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1083_out,
                 Y => SharedReg1084_out);

   SharedReg1085_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1084_out,
                 Y => SharedReg1085_out);

   SharedReg1086_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1085_out,
                 Y => SharedReg1086_out);

   SharedReg1087_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1086_out,
                 Y => SharedReg1087_out);

   SharedReg1088_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1087_out,
                 Y => SharedReg1088_out);

   SharedReg1089_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_8_impl_out,
                 Y => SharedReg1089_out);

   SharedReg1090_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1089_out,
                 Y => SharedReg1090_out);

   SharedReg1091_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1090_out,
                 Y => SharedReg1091_out);

   SharedReg1092_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1091_out,
                 Y => SharedReg1092_out);

   SharedReg1093_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1092_out,
                 Y => SharedReg1093_out);

   SharedReg1094_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1093_out,
                 Y => SharedReg1094_out);

   SharedReg1095_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1094_out,
                 Y => SharedReg1095_out);

   SharedReg1096_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1095_out,
                 Y => SharedReg1096_out);

   SharedReg1097_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1096_out,
                 Y => SharedReg1097_out);

   SharedReg1098_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1097_out,
                 Y => SharedReg1098_out);

   SharedReg1099_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1098_out,
                 Y => SharedReg1099_out);

   SharedReg1100_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1099_out,
                 Y => SharedReg1100_out);

   SharedReg1101_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1100_out,
                 Y => SharedReg1101_out);

   SharedReg1102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_0_impl_out,
                 Y => SharedReg1102_out);

   SharedReg1103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1102_out,
                 Y => SharedReg1103_out);

   SharedReg1104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1103_out,
                 Y => SharedReg1104_out);

   SharedReg1105_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1104_out,
                 Y => SharedReg1105_out);

   SharedReg1106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_1_impl_out,
                 Y => SharedReg1106_out);

   SharedReg1107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1106_out,
                 Y => SharedReg1107_out);

   SharedReg1108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1107_out,
                 Y => SharedReg1108_out);

   SharedReg1109_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1108_out,
                 Y => SharedReg1109_out);

   SharedReg1110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_0_impl_out,
                 Y => SharedReg1110_out);

   SharedReg1111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1110_out,
                 Y => SharedReg1111_out);

   SharedReg1112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1111_out,
                 Y => SharedReg1112_out);

   SharedReg1113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1112_out,
                 Y => SharedReg1113_out);

   SharedReg1114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1113_out,
                 Y => SharedReg1114_out);

   SharedReg1115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1114_out,
                 Y => SharedReg1115_out);

   SharedReg1116_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1115_out,
                 Y => SharedReg1116_out);

   SharedReg1117_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1116_out,
                 Y => SharedReg1117_out);

   SharedReg1118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_1_impl_out,
                 Y => SharedReg1118_out);

   SharedReg1119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1118_out,
                 Y => SharedReg1119_out);

   SharedReg1120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1119_out,
                 Y => SharedReg1120_out);

   SharedReg1121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1120_out,
                 Y => SharedReg1121_out);

   SharedReg1122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1121_out,
                 Y => SharedReg1122_out);

   SharedReg1123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1122_out,
                 Y => SharedReg1123_out);

   SharedReg1124_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1123_out,
                 Y => SharedReg1124_out);

   SharedReg1125_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1124_out,
                 Y => SharedReg1125_out);

   SharedReg1126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_2_impl_out,
                 Y => SharedReg1126_out);

   SharedReg1127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1126_out,
                 Y => SharedReg1127_out);

   SharedReg1128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1127_out,
                 Y => SharedReg1128_out);

   SharedReg1129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1128_out,
                 Y => SharedReg1129_out);

   SharedReg1130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1129_out,
                 Y => SharedReg1130_out);

   SharedReg1131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1130_out,
                 Y => SharedReg1131_out);

   SharedReg1132_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1131_out,
                 Y => SharedReg1132_out);

   SharedReg1133_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1132_out,
                 Y => SharedReg1133_out);

   SharedReg1134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_3_impl_out,
                 Y => SharedReg1134_out);

   SharedReg1135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1134_out,
                 Y => SharedReg1135_out);

   SharedReg1136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1135_out,
                 Y => SharedReg1136_out);

   SharedReg1137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1136_out,
                 Y => SharedReg1137_out);

   SharedReg1138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1137_out,
                 Y => SharedReg1138_out);

   SharedReg1139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1138_out,
                 Y => SharedReg1139_out);

   SharedReg1140_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1139_out,
                 Y => SharedReg1140_out);

   SharedReg1141_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1140_out,
                 Y => SharedReg1141_out);

   SharedReg1142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_4_impl_out,
                 Y => SharedReg1142_out);

   SharedReg1143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1142_out,
                 Y => SharedReg1143_out);

   SharedReg1144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1143_out,
                 Y => SharedReg1144_out);

   SharedReg1145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1144_out,
                 Y => SharedReg1145_out);

   SharedReg1146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1145_out,
                 Y => SharedReg1146_out);

   SharedReg1147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1146_out,
                 Y => SharedReg1147_out);

   SharedReg1148_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1147_out,
                 Y => SharedReg1148_out);

   SharedReg1149_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1148_out,
                 Y => SharedReg1149_out);

   SharedReg1150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_5_impl_out,
                 Y => SharedReg1150_out);

   SharedReg1151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1150_out,
                 Y => SharedReg1151_out);

   SharedReg1152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1151_out,
                 Y => SharedReg1152_out);

   SharedReg1153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1152_out,
                 Y => SharedReg1153_out);

   SharedReg1154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1153_out,
                 Y => SharedReg1154_out);

   SharedReg1155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1154_out,
                 Y => SharedReg1155_out);

   SharedReg1156_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1155_out,
                 Y => SharedReg1156_out);

   SharedReg1157_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1156_out,
                 Y => SharedReg1157_out);

   SharedReg1158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_6_impl_out,
                 Y => SharedReg1158_out);

   SharedReg1159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1158_out,
                 Y => SharedReg1159_out);

   SharedReg1160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1159_out,
                 Y => SharedReg1160_out);

   SharedReg1161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1160_out,
                 Y => SharedReg1161_out);

   SharedReg1162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1161_out,
                 Y => SharedReg1162_out);

   SharedReg1163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1162_out,
                 Y => SharedReg1163_out);

   SharedReg1164_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1163_out,
                 Y => SharedReg1164_out);

   SharedReg1165_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1164_out,
                 Y => SharedReg1165_out);

   SharedReg1166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_7_impl_out,
                 Y => SharedReg1166_out);

   SharedReg1167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1166_out,
                 Y => SharedReg1167_out);

   SharedReg1168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1167_out,
                 Y => SharedReg1168_out);

   SharedReg1169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1168_out,
                 Y => SharedReg1169_out);

   SharedReg1170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1169_out,
                 Y => SharedReg1170_out);

   SharedReg1171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1170_out,
                 Y => SharedReg1171_out);

   SharedReg1172_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1171_out,
                 Y => SharedReg1172_out);

   SharedReg1173_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1172_out,
                 Y => SharedReg1173_out);

   SharedReg1174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_8_impl_out,
                 Y => SharedReg1174_out);

   SharedReg1175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1174_out,
                 Y => SharedReg1175_out);

   SharedReg1176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1175_out,
                 Y => SharedReg1176_out);

   SharedReg1177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1176_out,
                 Y => SharedReg1177_out);

   SharedReg1178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1177_out,
                 Y => SharedReg1178_out);

   SharedReg1179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1178_out,
                 Y => SharedReg1179_out);

   SharedReg1180_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1179_out,
                 Y => SharedReg1180_out);

   SharedReg1181_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1180_out,
                 Y => SharedReg1181_out);

   SharedReg1182_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg1182_out);

   SharedReg1183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1182_out,
                 Y => SharedReg1183_out);

   SharedReg1184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1183_out,
                 Y => SharedReg1184_out);

   SharedReg1185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1184_out,
                 Y => SharedReg1185_out);

   SharedReg1186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1185_out,
                 Y => SharedReg1186_out);

   SharedReg1187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1186_out,
                 Y => SharedReg1187_out);

   SharedReg1188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1187_out,
                 Y => SharedReg1188_out);

   SharedReg1189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1188_out,
                 Y => SharedReg1189_out);

   SharedReg1190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1189_out,
                 Y => SharedReg1190_out);

   SharedReg1191_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1190_out,
                 Y => SharedReg1191_out);

   SharedReg1192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1191_out,
                 Y => SharedReg1192_out);

   SharedReg1193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1192_out,
                 Y => SharedReg1193_out);

   SharedReg1194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1193_out,
                 Y => SharedReg1194_out);

   SharedReg1195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1194_out,
                 Y => SharedReg1195_out);

   SharedReg1196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1195_out,
                 Y => SharedReg1196_out);

   SharedReg1197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1196_out,
                 Y => SharedReg1197_out);

   SharedReg1198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1197_out,
                 Y => SharedReg1198_out);

   SharedReg1199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1198_out,
                 Y => SharedReg1199_out);

   SharedReg1200_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1199_out,
                 Y => SharedReg1200_out);

   SharedReg1201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1200_out,
                 Y => SharedReg1201_out);

   SharedReg1202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1201_out,
                 Y => SharedReg1202_out);

   SharedReg1203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1202_out,
                 Y => SharedReg1203_out);

   SharedReg1204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1203_out,
                 Y => SharedReg1204_out);

   SharedReg1205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1204_out,
                 Y => SharedReg1205_out);

   SharedReg1206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1205_out,
                 Y => SharedReg1206_out);

   SharedReg1207_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1206_out,
                 Y => SharedReg1207_out);

   SharedReg1208_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1207_out,
                 Y => SharedReg1208_out);

   SharedReg1209_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1208_out,
                 Y => SharedReg1209_out);

   SharedReg1210_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg1210_out);

   SharedReg1211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1210_out,
                 Y => SharedReg1211_out);

   SharedReg1212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1211_out,
                 Y => SharedReg1212_out);

   SharedReg1213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1212_out,
                 Y => SharedReg1213_out);

   SharedReg1214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1213_out,
                 Y => SharedReg1214_out);

   SharedReg1215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1214_out,
                 Y => SharedReg1215_out);

   SharedReg1216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1215_out,
                 Y => SharedReg1216_out);

   SharedReg1217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1216_out,
                 Y => SharedReg1217_out);

   SharedReg1218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1217_out,
                 Y => SharedReg1218_out);

   SharedReg1219_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1218_out,
                 Y => SharedReg1219_out);

   SharedReg1220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1219_out,
                 Y => SharedReg1220_out);

   SharedReg1221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1220_out,
                 Y => SharedReg1221_out);

   SharedReg1222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1221_out,
                 Y => SharedReg1222_out);

   SharedReg1223_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1222_out,
                 Y => SharedReg1223_out);

   SharedReg1224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1223_out,
                 Y => SharedReg1224_out);

   SharedReg1225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1224_out,
                 Y => SharedReg1225_out);

   SharedReg1226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1225_out,
                 Y => SharedReg1226_out);

   SharedReg1227_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1226_out,
                 Y => SharedReg1227_out);

   SharedReg1228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1227_out,
                 Y => SharedReg1228_out);

   SharedReg1229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1228_out,
                 Y => SharedReg1229_out);

   SharedReg1230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1229_out,
                 Y => SharedReg1230_out);

   SharedReg1231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1230_out,
                 Y => SharedReg1231_out);

   SharedReg1232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1231_out,
                 Y => SharedReg1232_out);

   SharedReg1233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1232_out,
                 Y => SharedReg1233_out);

   SharedReg1234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1233_out,
                 Y => SharedReg1234_out);

   SharedReg1235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1234_out,
                 Y => SharedReg1235_out);

   SharedReg1236_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1235_out,
                 Y => SharedReg1236_out);

   SharedReg1237_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1236_out,
                 Y => SharedReg1237_out);

   SharedReg1238_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg1238_out);

   SharedReg1239_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1238_out,
                 Y => SharedReg1239_out);

   SharedReg1240_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1239_out,
                 Y => SharedReg1240_out);

   SharedReg1241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1240_out,
                 Y => SharedReg1241_out);

   SharedReg1242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1241_out,
                 Y => SharedReg1242_out);

   SharedReg1243_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg1243_out);

   SharedReg1244_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1243_out,
                 Y => SharedReg1244_out);

   SharedReg1245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1244_out,
                 Y => SharedReg1245_out);

   SharedReg1246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1245_out,
                 Y => SharedReg1246_out);

   SharedReg1247_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg1247_out);

   SharedReg1248_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg1248_out);

   SharedReg1249_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg1249_out);

   SharedReg1250_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1249_out,
                 Y => SharedReg1250_out);

   SharedReg1251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1250_out,
                 Y => SharedReg1251_out);

   SharedReg1252_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1251_out,
                 Y => SharedReg1252_out);

   SharedReg1253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1252_out,
                 Y => SharedReg1253_out);

   SharedReg1254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1253_out,
                 Y => SharedReg1254_out);

   SharedReg1255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1254_out,
                 Y => SharedReg1255_out);

   SharedReg1256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1255_out,
                 Y => SharedReg1256_out);

   SharedReg1257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1256_out,
                 Y => SharedReg1257_out);

   SharedReg1258_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg1258_out);

   SharedReg1259_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1258_out,
                 Y => SharedReg1259_out);

   SharedReg1260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1259_out,
                 Y => SharedReg1260_out);

   SharedReg1261_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1260_out,
                 Y => SharedReg1261_out);

   SharedReg1262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1261_out,
                 Y => SharedReg1262_out);

   SharedReg1263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1262_out,
                 Y => SharedReg1263_out);

   SharedReg1264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1263_out,
                 Y => SharedReg1264_out);

   SharedReg1265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1264_out,
                 Y => SharedReg1265_out);

   SharedReg1266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1265_out,
                 Y => SharedReg1266_out);

   SharedReg1267_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg1267_out);

   SharedReg1268_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1267_out,
                 Y => SharedReg1268_out);

   SharedReg1269_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg1269_out);

   SharedReg1270_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1269_out,
                 Y => SharedReg1270_out);

   SharedReg1271_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg1271_out);

   SharedReg1272_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1271_out,
                 Y => SharedReg1272_out);

   SharedReg1273_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1272_out,
                 Y => SharedReg1273_out);

   SharedReg1274_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1273_out,
                 Y => SharedReg1274_out);

   SharedReg1275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1274_out,
                 Y => SharedReg1275_out);

   SharedReg1276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1275_out,
                 Y => SharedReg1276_out);

   SharedReg1277_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg1277_out);

   SharedReg1278_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1277_out,
                 Y => SharedReg1278_out);

   SharedReg1279_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1278_out,
                 Y => SharedReg1279_out);

   SharedReg1280_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1279_out,
                 Y => SharedReg1280_out);

   SharedReg1281_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1280_out,
                 Y => SharedReg1281_out);

   SharedReg1282_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg1282_out);

   SharedReg1283_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1282_out,
                 Y => SharedReg1283_out);

   SharedReg1284_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg1284_out);

   SharedReg1285_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1284_out,
                 Y => SharedReg1285_out);

   SharedReg1286_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg1286_out);

   SharedReg1287_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg1287_out);

   SharedReg1288_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1287_out,
                 Y => SharedReg1288_out);
end architecture;

