--------------------------------------------------------------------------------
--                         ModuloCounter_3_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_3_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of ModuloCounter_3_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(1 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 2 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid3434711
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid3434711 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid3434711 is
signal XX_m3434712 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m3434712 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m3434712 <= X ;
   YY_m3434712 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid3434715
--                   (IntAdderClassical_33_f500_uid3434717)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid3434715 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid3434715 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid3434711 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid3434715 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid3434711  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid3434715  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_3_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_3_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_3_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid3435022_RightShifter
--                (RightShifter_24_by_max_26_F250_uid3435024)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid3435022_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid3435022_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid3435027
--                  (IntAdderAlternative_27_f250_uid3435031)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid3435027 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid3435027 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid3435034
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid3435034 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid3435034 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid3435037
--                   (IntAdderClassical_34_f250_uid3435039)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid3435037 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid3435037 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid3435022
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid3435022 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid3435022 is
   component FPAdd_8_23_uid3435022_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid3435027 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid3435034 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid3435037 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid3435022_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid3435027  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid3435034  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid3435037  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid3435022 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid3435022  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid3436309_RightShifter
--                (RightShifter_24_by_max_26_F250_uid3436311)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid3436309_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid3436309_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid3436314
--                  (IntAdderAlternative_27_f250_uid3436318)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid3436314 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid3436314 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid3436321
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid3436321 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid3436321 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid3436324
--                   (IntAdderClassical_34_f250_uid3436326)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid3436324 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid3436324 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid3436309
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid3436309 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid3436309 is
   component FPAdd_8_23_uid3436309_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid3436314 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid3436321 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid3436324 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid3436309_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid3436314  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid3436321  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid3436324  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid3436309 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid3436309  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 88 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      Y <= s87;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 90 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      Y <= s89;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 76 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      Y <= s75;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 95 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      Y <= s94;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 93 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      Y <= s92;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 87 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      Y <= s86;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 105 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      Y <= s104;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 82 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      Y <= s81;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 107 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      Y <= s106;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 62 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      Y <= s61;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 40 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      Y <= s39;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 71 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      Y <= s70;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "1" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 81 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      Y <= s80;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 74 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      Y <= s73;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1 : in std_logic_vector(31 downto 0);
          R_U : in std_logic_vector(31 downto 0);
          R_V : in std_logic_vector(31 downto 0);
          R_W : in std_logic_vector(31 downto 0);
          Inv_11 : out std_logic_vector(31 downto 0);
          Inv_12 : out std_logic_vector(31 downto 0);
          Inv_13 : out std_logic_vector(31 downto 0);
          Inv_21 : out std_logic_vector(31 downto 0);
          Inv_22 : out std_logic_vector(31 downto 0);
          Inv_23 : out std_logic_vector(31 downto 0);
          Inv_31 : out std_logic_vector(31 downto 0);
          Inv_32 : out std_logic_vector(31 downto 0);
          Inv_33 : out std_logic_vector(31 downto 0);
          Inv_41 : out std_logic_vector(31 downto 0);
          Inv_42 : out std_logic_vector(31 downto 0);
          Inv_43 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_3_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(1 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_3_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount31_out : std_logic_vector(1 downto 0) := (others => '0');
signal Ldiff_UU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add61_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product1010_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1010_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1010_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product101_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product101_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product101_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product121_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product121_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product141_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product141_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product161_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product161_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product161_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product171_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product171_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product171_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product181_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product191_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product191_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product191_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product241_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product271_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product271_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product271_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product331_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product331_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product351_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product351_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product351_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product411_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product412_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product412_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product412_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product58_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product58_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product58_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product59_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product60_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product60_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product60_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product64_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product65_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product65_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product65_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product66_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product72_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product74_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product74_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product74_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product76_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product77_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product77_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product77_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product81_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product81_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product81_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product84_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product84_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product84_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product86_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product86_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product86_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product87_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product87_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product87_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product88_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product88_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product88_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product94_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product94_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product94_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product97_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product97_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product97_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product98_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product98_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product98_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product99_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product99_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product99_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product34_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product40_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product40_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product43_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product43_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product44_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product44_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product47_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product47_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product49_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product49_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay23No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay47No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay31No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add24_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add61_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add61_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product74_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product74_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product76_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product76_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product77_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product77_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product81_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product81_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product84_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product84_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product86_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product86_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product87_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product87_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product88_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product88_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product94_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product94_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product97_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product97_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product98_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product98_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product99_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product99_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract3_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract3_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add112_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add112_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add12_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add12_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add15_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add15_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add4_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add4_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add7_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add7_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add9_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add9_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product116_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product116_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product10_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product10_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product13_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product13_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product16_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product16_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product18_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product18_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product19_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product19_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product21_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product21_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product23_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product23_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product28_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product28_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product31_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product31_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product34_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product34_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product4_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product4_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product40_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product40_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product43_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product43_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product44_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product44_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product47_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product47_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product49_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product49_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product6_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product6_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay93No1_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No1_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No1_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No2_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add110_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add110_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No35_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add101_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add101_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No7_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No7_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add121_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add121_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add131_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add131_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No13_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay23No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No3_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay31No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No2_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add61_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add61_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product1010_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product1010_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product101_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product101_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product114_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product114_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product121_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product121_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product141_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product141_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product161_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product161_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product171_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product171_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product181_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product181_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product191_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product191_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No1_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product241_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product241_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product271_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product271_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product312_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product312_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product321_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product321_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product331_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product331_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product351_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product351_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product411_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product411_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No38_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product412_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product412_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product512_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product512_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product58_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product58_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product59_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product59_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product60_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product60_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product64_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product64_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product65_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product65_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No42_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product66_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product66_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product72_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product72_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product74_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product74_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product76_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product76_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product77_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product77_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product81_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product81_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product84_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product84_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No2_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product86_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product86_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product87_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product87_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No11_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product88_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product88_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product94_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product94_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product97_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product97_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product98_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product98_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product99_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product99_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No3_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No5_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay47No_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Add112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Add112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No1_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Add12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Add12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay63No_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Add15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Add15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay33No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Add4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Add4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay30No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Add7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Add7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay35No_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Add9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Add9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Divide_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Divide_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product10_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product10_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No15_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product28_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product28_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product31_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product31_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product34_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product34_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product40_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product40_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product43_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product43_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product44_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product44_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product47_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product47_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product49_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product49_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount31_instance: ModuloCounter_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount31_out);
Ldiff_UU_del_1_IEEE <= Ldiff_UU_del_1;
   Ldiff_UU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_out,
                 X => Ldiff_UU_del_1_IEEE);
Ldiff_UV_del_1_IEEE <= Ldiff_UV_del_1;
   Ldiff_UV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_out,
                 X => Ldiff_UV_del_1_IEEE);
Ldiff_UW_del_1_IEEE <= Ldiff_UW_del_1;
   Ldiff_UW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_out,
                 X => Ldiff_UW_del_1_IEEE);
Ldiff_VU_del_1_IEEE <= Ldiff_VU_del_1;
   Ldiff_VU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_out,
                 X => Ldiff_VU_del_1_IEEE);
Ldiff_VV_del_1_IEEE <= Ldiff_VV_del_1;
   Ldiff_VV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_out,
                 X => Ldiff_VV_del_1_IEEE);
Ldiff_VW_del_1_IEEE <= Ldiff_VW_del_1;
   Ldiff_VW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_out,
                 X => Ldiff_VW_del_1_IEEE);
Ldiff_WU_del_1_IEEE <= Ldiff_WU_del_1;
   Ldiff_WU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_out,
                 X => Ldiff_WU_del_1_IEEE);
Ldiff_WV_del_1_IEEE <= Ldiff_WV_del_1;
   Ldiff_WV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_out,
                 X => Ldiff_WV_del_1_IEEE);
Ldiff_WW_del_1_IEEE <= Ldiff_WW_del_1;
   Ldiff_WW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_out,
                 X => Ldiff_WW_del_1_IEEE);
R_U_IEEE <= R_U;
   R_U_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_out,
                 X => R_U_IEEE);
R_V_IEEE <= R_V;
   R_V_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_out,
                 X => R_V_IEEE);
R_W_IEEE <= R_W;
   R_W_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_out,
                 X => R_W_IEEE);

Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_impl_out,
                 X => Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg154_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg75_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_3_cast <= SharedReg75_out;
   MUX_Product108_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product108_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_impl_0_out,
                 Y => Delay1No_out);

SharedReg176_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
Delay90No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast <= Delay90No_out;
SharedReg17_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
   MUX_Product108_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay90No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product108_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product110_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_impl_out,
                 X => Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast);

SharedReg135_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg154_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg1_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
   MUX_Product110_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product110_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_impl_0_out,
                 Y => Delay1No2_out);

SharedReg183_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
Delay97No_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast <= Delay97No_out;
SharedReg16_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
   MUX_Product110_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product110_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product109_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_impl_out,
                 X => Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg154_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg93_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_3_cast <= SharedReg93_out;
   MUX_Product109_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg93_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product109_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_impl_0_out,
                 Y => Delay1No4_out);

SharedReg183_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg59_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast <= SharedReg59_out;
SharedReg185_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_3_cast <= SharedReg185_out;
   MUX_Product109_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg185_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product109_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product111_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_impl_out,
                 X => Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast);

SharedReg34_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg154_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg78_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast <= SharedReg78_out;
   MUX_Product111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg78_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product111_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_0_out,
                 Y => Delay1No6_out);

SharedReg178_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg178_out;
Delay79No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast <= Delay79No_out;
SharedReg175_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
   MUX_Product111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay79No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product111_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product210_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_impl_out,
                 X => Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast);

Delay7No2_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast <= Delay7No2_out;
SharedReg154_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg82_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
   MUX_Product210_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No2_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg82_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product210_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_0_out,
                 Y => Delay1No8_out);

SharedReg153_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
Delay97No1_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast <= Delay97No1_out;
SharedReg7_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast <= SharedReg7_out;
   MUX_Product210_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No1_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg7_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product210_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product310_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_impl_out,
                 X => Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg154_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg174_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product310_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product310_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_0_out,
                 Y => Delay1No10_out);

SharedReg29_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
Delay94No_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast <= Delay94No_out;
SharedReg174_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product310_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay94No_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product310_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product410_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_impl_out,
                 X => Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg154_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg87_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_3_cast <= SharedReg87_out;
   MUX_Product410_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg87_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product410_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_impl_0_out,
                 Y => Delay1No12_out);

SharedReg3_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast <= SharedReg3_out;
Delay89No_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast <= Delay89No_out;
SharedReg150_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
   MUX_Product410_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay89No_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product410_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product510_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_impl_out,
                 X => Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast);

SharedReg41_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg154_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg90_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
   MUX_Product510_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product510_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_impl_0_out,
                 Y => Delay1No14_out);

SharedReg29_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
Delay93No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast <= Delay93No_out;
SharedReg17_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
   MUX_Product510_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay93No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product510_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product610_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_impl_out,
                 X => Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast);

SharedReg77_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast <= SharedReg77_out;
SharedReg154_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg92_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_3_cast <= SharedReg92_out;
   MUX_Product610_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg77_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg92_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product610_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_impl_0_out,
                 Y => Delay1No16_out);

SharedReg148_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast <= SharedReg148_out;
Delay93No1_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast <= Delay93No1_out;
SharedReg7_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_3_cast <= SharedReg7_out;
   MUX_Product610_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay93No1_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg7_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product610_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product710_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_impl_out,
                 X => Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast);

Delay8No1_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast <= Delay8No1_out;
SharedReg154_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg174_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product710_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No1_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product710_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_impl_0_out,
                 Y => Delay1No18_out);

SharedReg153_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg55_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast <= SharedReg55_out;
SharedReg174_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product710_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product710_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product810_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_impl_out,
                 X => Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast);

SharedReg107_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg154_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg174_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product810_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product810_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_impl_0_out,
                 Y => Delay1No20_out);

SharedReg18_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg56_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast <= SharedReg56_out;
SharedReg174_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product810_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg56_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product810_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product910_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_impl_out,
                 X => Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast);

SharedReg86_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg154_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg94_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
   MUX_Product910_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product910_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_impl_0_out,
                 Y => Delay1No22_out);

SharedReg8_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg71_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg12_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_3_cast <= SharedReg12_out;
   MUX_Product910_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg12_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product910_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_impl_1_out,
                 Y => Delay1No23_out);
   Inv_11_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_IEEE,
                 X => Delay1No24_out);
Inv_11 <= Inv_11_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => Delay1No24_out);
   Inv_12_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_IEEE,
                 X => Delay1No25_out);
Inv_12 <= Inv_12_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => Delay1No25_out);
   Inv_13_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_IEEE,
                 X => Delay1No26_out);
Inv_13 <= Inv_13_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => Delay1No26_out);
   Inv_21_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_IEEE,
                 X => Delay1No27_out);
Inv_21 <= Inv_21_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => Delay1No27_out);
   Inv_22_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_IEEE,
                 X => Delay1No28_out);
Inv_22 <= Inv_22_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => Delay1No28_out);
   Inv_23_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_IEEE,
                 X => Delay1No29_out);
Inv_23 <= Inv_23_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay1No29_out);
   Inv_31_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_IEEE,
                 X => Delay1No30_out);
Inv_31 <= Inv_31_IEEE;

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => Delay1No30_out);
   Inv_32_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_IEEE,
                 X => Delay1No31_out);
Inv_32 <= Inv_32_IEEE;

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => Delay1No31_out);
   Inv_33_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_IEEE,
                 X => Delay1No32_out);
Inv_33 <= Inv_33_IEEE;

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => Delay1No32_out);
   Inv_41_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_IEEE,
                 X => Delay1No33_out);
Inv_41 <= Inv_41_IEEE;

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => Delay1No33_out);
   Inv_42_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_IEEE,
                 X => Delay1No34_out);
Inv_42 <= Inv_42_IEEE;

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => Delay1No34_out);
   Inv_43_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_IEEE,
                 X => Delay1No35_out);
Inv_43 <= Inv_43_IEEE;

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add30_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_impl_out,
                 X => Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
Delay89No1_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast <= Delay89No1_out;
SharedReg110_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_3_cast <= SharedReg110_out;
   MUX_Add30_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay89No1_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg110_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add30_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_impl_0_out,
                 Y => Delay1No36_out);

SharedReg119_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast <= SharedReg119_out;
Delay89No2_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast <= Delay89No2_out;
SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_3_cast <= SharedReg112_out;
   MUX_Add30_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg119_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay89No2_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add30_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add110_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add110_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add110_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_impl_out,
                 X => Delay1No38_out_to_Add110_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add110_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
Delay107No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast <= Delay107No_out;
Delay103No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_3_cast <= Delay103No_out;
   MUX_Add110_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay107No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay103No_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add110_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_impl_0_out,
                 Y => Delay1No38_out);

Delay2No35_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast <= Delay2No35_out;
SharedReg141_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
Delay96No_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_3_cast <= Delay96No_out;
   MUX_Add110_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No35_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay96No_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add110_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add101_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add101_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add101_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_impl_out,
                 X => Delay1No40_out_to_Add101_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add101_impl_parent_implementedSystem_port_1_cast);

SharedReg52_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg40_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg89_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_3_cast <= SharedReg89_out;
   MUX_Add101_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg89_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add101_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_impl_0_out,
                 Y => Delay1No40_out);

Delay3No7_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast <= Delay3No7_out;
SharedReg41_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg72_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_3_cast <= SharedReg72_out;
   MUX_Add101_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No7_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg72_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add101_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add111_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add111_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add111_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_impl_out,
                 X => Delay1No42_out_to_Add111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add111_impl_parent_implementedSystem_port_1_cast);

Delay10No7_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast <= Delay10No7_out;
SharedReg42_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg42_out;
Delay15No2_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast <= Delay15No2_out;
   MUX_Add111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay10No7_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay15No2_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add111_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_0_out,
                 Y => Delay1No42_out);

SharedReg139_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg139_out;
SharedReg44_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg44_out;
SharedReg73_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast <= SharedReg73_out;
   MUX_Add111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg139_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg44_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg73_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add111_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add121_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add121_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add121_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_impl_out,
                 X => Delay1No44_out_to_Add121_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add121_impl_parent_implementedSystem_port_1_cast);

SharedReg79_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast <= SharedReg79_out;
Delay20No_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast <= Delay20No_out;
SharedReg38_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast <= SharedReg38_out;
   MUX_Add121_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay20No_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg38_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add121_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_impl_0_out,
                 Y => Delay1No44_out);

SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast <= SharedReg102_out;
SharedReg137_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast <= SharedReg137_out;
Delay6No10_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast <= Delay6No10_out;
   MUX_Add121_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay6No10_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add121_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add131_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add131_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add131_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_impl_out,
                 X => Delay1No46_out_to_Add131_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add131_impl_parent_implementedSystem_port_1_cast);

SharedReg100_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg119_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast <= SharedReg119_out;
SharedReg36_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_3_cast <= SharedReg36_out;
   MUX_Add131_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add131_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_0_out,
                 Y => Delay1No46_out);

Delay3No13_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast <= Delay3No13_out;
SharedReg168_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast <= SharedReg168_out;
SharedReg61_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_3_cast <= SharedReg61_out;
   MUX_Add131_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No13_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg168_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg61_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add131_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add18_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_impl_out,
                 X => Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast);

SharedReg127_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
Delay61No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast <= Delay61No_out;
Delay23No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast <= Delay23No_out;
   MUX_Add18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay61No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay23No_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add18_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_0_out,
                 Y => Delay1No48_out);

SharedReg128_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg128_out;
SharedReg74_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg74_out;
SharedReg140_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast <= SharedReg140_out;
   MUX_Add18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg128_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg74_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg140_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add18_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add19_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add19_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add19_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add19_impl_out,
                 X => Delay1No50_out_to_Add19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add19_impl_parent_implementedSystem_port_1_cast);

Delay14No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast <= Delay14No_out;
SharedReg117_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
Delay18No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_3_cast <= Delay18No_out;
   MUX_Add19_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay14No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay18No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add19_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_impl_0_out,
                 Y => Delay1No50_out);

SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg143_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast <= SharedReg143_out;
SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
   MUX_Add19_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg143_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg65_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add19_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add20_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add20_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add20_impl_out,
                 X => Delay1No52_out_to_Add20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add20_impl_parent_implementedSystem_port_1_cast);

Delay18No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast <= Delay18No1_out;
Delay25No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast <= Delay25No1_out;
Delay11No3_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_3_cast <= Delay11No3_out;
   MUX_Add20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay18No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay25No1_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay11No3_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add20_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_0_out,
                 Y => Delay1No52_out);

SharedReg140_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg140_out;
SharedReg144_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg144_out;
SharedReg138_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_3_cast <= SharedReg138_out;
   MUX_Add20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg140_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg144_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg138_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add20_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add21_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add21_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add21_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add21_impl_out,
                 X => Delay1No54_out_to_Add21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add21_impl_parent_implementedSystem_port_1_cast);

SharedReg98_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg98_out;
Delay31No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast <= Delay31No_out;
Delay12No2_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_3_cast <= Delay12No2_out;
   MUX_Add21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay31No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay12No2_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add21_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_impl_0_out,
                 Y => Delay1No54_out);

SharedReg69_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg145_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
SharedReg141_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_3_cast <= SharedReg141_out;
   MUX_Add21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg141_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add21_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add22_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add22_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add22_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add22_impl_out,
                 X => Delay1No56_out_to_Add22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add22_impl_parent_implementedSystem_port_1_cast);

SharedReg133_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast <= SharedReg133_out;
Delay44No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast <= Delay44No_out;
Delay15No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast <= Delay15No_out;
   MUX_Add22_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay44No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay15No_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add22_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_0_out,
                 Y => Delay1No56_out);

SharedReg91_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast <= SharedReg142_out;
SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
   MUX_Add22_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Add22_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add24_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add24_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add24_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_impl_out,
                 X => Delay1No58_out_to_Add24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add24_impl_parent_implementedSystem_port_1_cast);

SharedReg46_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast <= SharedReg46_out;
Delay12No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast <= Delay12No4_out;
   MUX_Add24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay12No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add24_impl_0_LUT_out,
                 oMux => MUX_Add24_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_0_out,
                 Y => Delay1No58_out);

SharedReg48_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg137_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast <= SharedReg137_out;
   MUX_Add24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add24_impl_1_LUT_out,
                 oMux => MUX_Add24_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add61_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add61_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add61_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add61_impl_out,
                 X => Delay1No60_out_to_Add61_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add61_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
Delay65No_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast <= Delay65No_out;
   MUX_Add61_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay65No_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add61_impl_0_LUT_out,
                 oMux => MUX_Add61_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_0_out,
                 Y => Delay1No60_out);

SharedReg97_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg151_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
   MUX_Add61_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add61_impl_1_LUT_out,
                 oMux => MUX_Add61_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product112_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product112_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product112_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_impl_out,
                 X => Delay1No62_out_to_Product112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product112_impl_parent_implementedSystem_port_1_cast);

SharedReg124_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg173_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg50_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_3_cast <= SharedReg50_out;
   MUX_Product112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg50_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product112_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_0_out,
                 Y => Delay1No62_out);

SharedReg183_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg173_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg19_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
   MUX_Product112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg19_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product112_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product1010_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product1010_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product1010_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product1010_impl_out,
                 X => Delay1No64_out_to_Product1010_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product1010_impl_parent_implementedSystem_port_1_cast);

SharedReg94_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg173_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product1010_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product1010_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product1010_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1010_impl_0_out,
                 Y => Delay1No64_out);

SharedReg23_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg173_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product1010_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product1010_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product1010_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1010_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product101_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product101_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product101_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product101_impl_out,
                 X => Delay1No66_out_to_Product101_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product101_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg99_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_3_cast <= SharedReg99_out;
   MUX_Product101_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg99_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product101_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product101_impl_0_out,
                 Y => Delay1No66_out);

SharedReg13_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg7_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_3_cast <= SharedReg7_out;
   MUX_Product101_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg7_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product101_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product101_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product114_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product114_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product114_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_impl_out,
                 X => Delay1No68_out_to_Product114_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product114_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg76_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast <= SharedReg76_out;
SharedReg174_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product114_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product114_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_impl_0_out,
                 Y => Delay1No68_out);

SharedReg13_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg151_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
SharedReg174_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product114_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product114_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product121_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product121_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product121_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product121_impl_out,
                 X => Delay1No70_out_to_Product121_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product121_impl_parent_implementedSystem_port_1_cast);

SharedReg125_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg173_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg101_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_3_cast <= SharedReg101_out;
   MUX_Product121_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg101_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product121_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product121_impl_0_out,
                 Y => Delay1No70_out);

SharedReg176_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg22_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
   MUX_Product121_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg22_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product121_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product121_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product141_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product141_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product141_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product141_impl_out,
                 X => Delay1No72_out_to_Product141_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product141_impl_parent_implementedSystem_port_1_cast);

SharedReg126_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast <= SharedReg126_out;
SharedReg173_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product141_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg126_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product141_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product141_impl_0_out,
                 Y => Delay1No72_out);

SharedReg3_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg173_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product141_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product141_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product141_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product161_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product161_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product161_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product161_impl_out,
                 X => Delay1No74_out_to_Product161_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product161_impl_parent_implementedSystem_port_1_cast);

SharedReg129_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_1_cast <= SharedReg129_out;
SharedReg173_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product161_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg129_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product161_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product161_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product161_impl_0_out,
                 Y => Delay1No74_out);

SharedReg183_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg173_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product161_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product161_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product161_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product161_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product171_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product171_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product171_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product171_impl_out,
                 X => Delay1No76_out_to_Product171_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product171_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg173_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product171_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product171_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product171_impl_0_out,
                 Y => Delay1No76_out);

SharedReg183_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg173_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product171_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product171_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product171_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product181_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product181_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product181_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product181_impl_out,
                 X => Delay1No78_out_to_Product181_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product181_impl_parent_implementedSystem_port_1_cast);

SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg173_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg85_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_3_cast <= SharedReg85_out;
   MUX_Product181_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg85_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product181_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_impl_0_out,
                 Y => Delay1No78_out);

SharedReg176_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg147_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_3_cast <= SharedReg147_out;
   MUX_Product181_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg147_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product181_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product191_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product191_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product191_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product191_impl_out,
                 X => Delay1No80_out_to_Product191_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product191_impl_parent_implementedSystem_port_1_cast);

SharedReg148_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg173_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product191_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product191_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product191_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product191_impl_0_out,
                 Y => Delay1No80_out);

Delay12No1_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_1_cast <= Delay12No1_out;
SharedReg173_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product191_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No1_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product191_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product191_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product191_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product241_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product241_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product241_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product241_impl_out,
                 X => Delay1No82_out_to_Product241_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product241_impl_parent_implementedSystem_port_1_cast);

SharedReg156_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast <= SharedReg156_out;
SharedReg173_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product241_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg156_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product241_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_0_out,
                 Y => Delay1No82_out);

Delay21No_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast <= Delay21No_out;
SharedReg173_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product241_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay21No_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product241_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product271_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product271_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product271_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product271_impl_out,
                 X => Delay1No84_out_to_Product271_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product271_impl_parent_implementedSystem_port_1_cast);

SharedReg157_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast <= SharedReg157_out;
SharedReg173_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
Delay7No4_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_3_cast <= Delay7No4_out;
   MUX_Product271_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg157_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay7No4_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product271_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product271_impl_0_out,
                 Y => Delay1No84_out);

SharedReg186_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg173_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg150_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
   MUX_Product271_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product271_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product271_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product312_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product312_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product312_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_impl_out,
                 X => Delay1No86_out_to_Product312_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product312_impl_parent_implementedSystem_port_1_cast);

SharedReg158_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast <= SharedReg158_out;
SharedReg96_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast <= SharedReg96_out;
SharedReg124_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_3_cast <= SharedReg124_out;
   MUX_Product312_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg158_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg96_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg124_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product312_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_0_out,
                 Y => Delay1No86_out);

SharedReg178_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg24_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg182_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_3_cast <= SharedReg182_out;
   MUX_Product312_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg182_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product312_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product321_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product321_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product321_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_impl_out,
                 X => Delay1No88_out_to_Product321_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product321_impl_parent_implementedSystem_port_1_cast);

SharedReg155_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast <= SharedReg155_out;
SharedReg173_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
Delay6No12_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast <= Delay6No12_out;
   MUX_Product321_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg155_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay6No12_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product321_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_0_out,
                 Y => Delay1No88_out);

SharedReg186_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg173_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg150_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
   MUX_Product321_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product321_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product331_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product331_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product331_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product331_impl_out,
                 X => Delay1No90_out_to_Product331_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product331_impl_parent_implementedSystem_port_1_cast);

SharedReg160_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg173_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg109_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_3_cast <= SharedReg109_out;
   MUX_Product331_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg109_out_to_MUX_Product331_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product331_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_impl_0_out,
                 Y => Delay1No90_out);

SharedReg186_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg173_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg28_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
   MUX_Product331_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg28_out_to_MUX_Product331_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product331_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product331_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product351_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product351_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product351_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product351_impl_out,
                 X => Delay1No92_out_to_Product351_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product351_impl_parent_implementedSystem_port_1_cast);

Delay2No36_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_1_cast <= Delay2No36_out;
SharedReg173_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product351_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No36_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product351_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product351_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product351_impl_0_out,
                 Y => Delay1No92_out);

SharedReg183_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg173_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product351_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product351_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product351_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product351_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product411_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product411_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product411_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product411_impl_out,
                 X => Delay1No94_out_to_Product411_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product411_impl_parent_implementedSystem_port_1_cast);

Delay2No38_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_1_cast <= Delay2No38_out;
SharedReg173_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product411_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No38_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product411_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product411_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_impl_0_out,
                 Y => Delay1No94_out);

SharedReg176_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product411_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product411_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product411_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product412_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product412_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product412_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product412_impl_out,
                 X => Delay1No96_out_to_Product412_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product412_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg173_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg111_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_3_cast <= SharedReg111_out;
   MUX_Product412_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product412_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product412_impl_0_out,
                 Y => Delay1No96_out);

SharedReg181_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg173_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg28_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
   MUX_Product412_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg28_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product412_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product412_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product512_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product512_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product512_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_impl_out,
                 X => Delay1No98_out_to_Product512_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product512_impl_parent_implementedSystem_port_1_cast);

SharedReg164_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg173_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg113_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_3_cast <= SharedReg113_out;
   MUX_Product512_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg113_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product512_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_impl_0_out,
                 Y => Delay1No98_out);

SharedReg186_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg173_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg2_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
   MUX_Product512_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product512_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product57_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product57_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product57_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product57_impl_out,
                 X => Delay1No100_out_to_Product57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product57_impl_parent_implementedSystem_port_1_cast);

SharedReg161_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg173_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg115_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
   MUX_Product57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product57_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_impl_0_out,
                 Y => Delay1No100_out);

SharedReg178_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg173_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg22_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
   MUX_Product57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg22_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product57_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product58_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product58_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product58_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product58_impl_out,
                 X => Delay1No102_out_to_Product58_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product58_impl_parent_implementedSystem_port_1_cast);

SharedReg167_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_1_cast <= SharedReg167_out;
SharedReg173_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product58_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product58_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product58_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product58_impl_0_out,
                 Y => Delay1No102_out);

SharedReg178_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg173_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg174_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
   MUX_Product58_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product58_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product58_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product58_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product59_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product59_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product59_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product59_impl_out,
                 X => Delay1No104_out_to_Product59_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product59_impl_parent_implementedSystem_port_1_cast);

SharedReg165_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg173_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg119_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_3_cast <= SharedReg119_out;
   MUX_Product59_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg119_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product59_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_impl_0_out,
                 Y => Delay1No104_out);

SharedReg176_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg2_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
   MUX_Product59_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product59_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product60_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product60_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product60_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product60_impl_out,
                 X => Delay1No106_out_to_Product60_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product60_impl_parent_implementedSystem_port_1_cast);

SharedReg166_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg104_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg120_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_3_cast <= SharedReg120_out;
   MUX_Product60_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product60_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product60_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product60_impl_0_out,
                 Y => Delay1No106_out);

SharedReg186_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg146_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
SharedReg12_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_3_cast <= SharedReg12_out;
   MUX_Product60_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg12_out_to_MUX_Product60_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product60_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product60_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product64_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product64_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product64_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product64_impl_out,
                 X => Delay1No108_out_to_Product64_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product64_impl_parent_implementedSystem_port_1_cast);

SharedReg171_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg173_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg106_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_3_cast <= SharedReg106_out;
   MUX_Product64_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg106_out_to_MUX_Product64_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product64_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_impl_0_out,
                 Y => Delay1No108_out);

SharedReg186_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg173_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg152_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_3_cast <= SharedReg152_out;
   MUX_Product64_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg152_out_to_MUX_Product64_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product64_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product65_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product65_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product65_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product65_impl_out,
                 X => Delay1No110_out_to_Product65_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product65_impl_parent_implementedSystem_port_1_cast);

Delay2No42_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast <= Delay2No42_out;
SharedReg173_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg123_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_3_cast <= SharedReg123_out;
   MUX_Product65_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No42_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg123_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product65_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product65_impl_0_out,
                 Y => Delay1No110_out);

SharedReg176_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg147_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_3_cast <= SharedReg147_out;
   MUX_Product65_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg147_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product65_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product65_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product66_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product66_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product66_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product66_impl_out,
                 X => Delay1No112_out_to_Product66_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product66_impl_parent_implementedSystem_port_1_cast);

SharedReg172_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast <= SharedReg172_out;
SharedReg173_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg114_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_3_cast <= SharedReg114_out;
   MUX_Product66_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg172_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg114_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product66_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_impl_0_out,
                 Y => Delay1No112_out);

SharedReg176_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg173_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
SharedReg150_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
   MUX_Product66_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product66_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product72_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product72_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product72_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product72_impl_out,
                 X => Delay1No114_out_to_Product72_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product72_impl_parent_implementedSystem_port_1_cast);

Delay12No_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast <= Delay12No_out;
SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg150_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_3_cast <= SharedReg150_out;
   MUX_Product72_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product72_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_0_out,
                 Y => Delay1No114_out);

SharedReg153_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg151_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
Delay11No1_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_3_cast <= Delay11No1_out;
   MUX_Product72_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay11No1_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Product72_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product74_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product74_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product74_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product74_impl_out,
                 X => Delay1No116_out_to_Product74_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product74_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg15_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product74_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product74_impl_0_LUT_out,
                 oMux => MUX_Product74_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product74_impl_0_out,
                 Y => Delay1No116_out);

SharedReg26_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Product74_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product74_impl_1_LUT_out,
                 oMux => MUX_Product74_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product74_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product76_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product76_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product76_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product76_impl_out,
                 X => Delay1No118_out_to_Product76_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product76_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg174_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
   MUX_Product76_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product76_impl_0_LUT_out,
                 oMux => MUX_Product76_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_impl_0_out,
                 Y => Delay1No118_out);

SharedReg151_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg174_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast <= SharedReg174_out;
   MUX_Product76_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product76_impl_1_LUT_out,
                 oMux => MUX_Product76_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product77_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product77_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product77_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product77_impl_out,
                 X => Delay1No120_out_to_Product77_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product77_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg126_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast <= SharedReg126_out;
   MUX_Product77_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product77_impl_0_LUT_out,
                 oMux => MUX_Product77_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product77_impl_0_out,
                 Y => Delay1No120_out);

SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg182_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product77_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product77_impl_1_LUT_out,
                 oMux => MUX_Product77_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product77_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product81_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product81_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product81_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product81_impl_out,
                 X => Delay1No122_out_to_Product81_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product81_impl_parent_implementedSystem_port_1_cast);

SharedReg125_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg127_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast <= SharedReg127_out;
   MUX_Product81_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product81_impl_0_LUT_out,
                 oMux => MUX_Product81_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product81_impl_0_out,
                 Y => Delay1No122_out);

SharedReg177_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg175_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Product81_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product81_impl_1_LUT_out,
                 oMux => MUX_Product81_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product81_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product84_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product84_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product84_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product84_impl_out,
                 X => Delay1No124_out_to_Product84_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product84_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg147_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast <= SharedReg147_out;
   MUX_Product84_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product84_impl_0_LUT_out,
                 oMux => MUX_Product84_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product84_impl_0_out,
                 Y => Delay1No124_out);

Delay11No2_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast <= Delay11No2_out;
SharedReg151_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
   MUX_Product84_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No2_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product84_impl_1_LUT_out,
                 oMux => MUX_Product84_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product84_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product86_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product86_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product86_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product86_impl_out,
                 X => Delay1No126_out_to_Product86_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product86_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg6_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
   MUX_Product86_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Product86_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product86_impl_0_LUT_out,
                 oMux => MUX_Product86_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product86_impl_0_out,
                 Y => Delay1No126_out);

SharedReg21_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Product86_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product86_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product86_impl_1_LUT_out,
                 oMux => MUX_Product86_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product86_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product87_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product87_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product87_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product87_impl_out,
                 X => Delay1No128_out_to_Product87_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product87_impl_parent_implementedSystem_port_1_cast);

Delay3No11_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast <= Delay3No11_out;
SharedReg146_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product87_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No11_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product87_impl_0_LUT_out,
                 oMux => MUX_Product87_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product87_impl_0_out,
                 Y => Delay1No128_out);

SharedReg151_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg185_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast <= SharedReg185_out;
   MUX_Product87_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product87_impl_1_LUT_out,
                 oMux => MUX_Product87_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product87_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product88_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product88_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product88_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product88_impl_out,
                 X => Delay1No130_out_to_Product88_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product88_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg130_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product88_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product88_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product88_impl_0_LUT_out,
                 oMux => MUX_Product88_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product88_impl_0_out,
                 Y => Delay1No130_out);

SharedReg21_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg175_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Product88_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product88_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product88_impl_1_LUT_out,
                 oMux => MUX_Product88_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product88_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product94_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product94_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product94_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product94_impl_out,
                 X => Delay1No132_out_to_Product94_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product94_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg132_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product94_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product94_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product94_impl_0_LUT_out,
                 oMux => MUX_Product94_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product94_impl_0_out,
                 Y => Delay1No132_out);

SharedReg21_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg180_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_2_cast <= SharedReg180_out;
   MUX_Product94_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg180_out_to_MUX_Product94_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product94_impl_1_LUT_out,
                 oMux => MUX_Product94_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product94_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product97_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product97_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product97_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product97_impl_out,
                 X => Delay1No134_out_to_Product97_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product97_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg146_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product97_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product97_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product97_impl_0_LUT_out,
                 oMux => MUX_Product97_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product97_impl_0_out,
                 Y => Delay1No134_out);

SharedReg11_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg20_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
   MUX_Product97_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product97_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product97_impl_1_LUT_out,
                 oMux => MUX_Product97_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product97_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product98_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product98_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product98_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product98_impl_out,
                 X => Delay1No136_out_to_Product98_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product98_impl_parent_implementedSystem_port_1_cast);

Delay11No_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast <= Delay11No_out;
SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
   MUX_Product98_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product98_impl_0_LUT_out,
                 oMux => MUX_Product98_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product98_impl_0_out,
                 Y => Delay1No136_out);

SharedReg150_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg149_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast <= SharedReg149_out;
   MUX_Product98_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product98_impl_1_LUT_out,
                 oMux => MUX_Product98_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product98_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product99_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product99_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product99_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product99_impl_out,
                 X => Delay1No138_out_to_Product99_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product99_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg147_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast <= SharedReg147_out;
   MUX_Product99_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product99_impl_0_LUT_out,
                 oMux => MUX_Product99_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product99_impl_0_out,
                 Y => Delay1No138_out);

SharedReg21_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg150_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast <= SharedReg150_out;
   MUX_Product99_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg150_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product99_impl_1_LUT_out,
                 oMux => MUX_Product99_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product99_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Subtract12_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_impl_out,
                 X => Delay1No140_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast);

Delay12No3_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast <= Delay12No3_out;
Delay17No_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast <= Delay17No_out;
SharedReg83_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_3_cast <= SharedReg83_out;
   MUX_Subtract12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No3_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay17No_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg83_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract12_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_0_out,
                 Y => Delay1No140_out);

SharedReg54_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg57_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg57_out;
Delay2No17_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_3_cast <= Delay2No17_out;
   MUX_Subtract12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No17_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract12_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract1_impl_out,
                 X => Delay1No142_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg108_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg108_out;
Delay8No2_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_3_cast <= Delay8No2_out;
   MUX_Subtract1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay8No2_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract1_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_impl_0_out,
                 Y => Delay1No142_out);

SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg53_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
   MUX_Subtract1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract1_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Subtract11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract11_impl_out,
                 X => Delay1No144_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast);

Delay9No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast <= Delay9No_out;
Delay22No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast <= Delay22No_out;
Delay8No3_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast <= Delay8No3_out;
   MUX_Subtract11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay9No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay22No_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay8No3_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract11_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_0_out,
                 Y => Delay1No144_out);

SharedReg63_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg67_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg67_out;
SharedReg60_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast <= SharedReg60_out;
   MUX_Subtract11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg67_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg60_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => ModCount31_out,
                 oMux => MUX_Subtract11_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Subtract2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_impl_out,
                 X => Delay1No146_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast);

SharedReg42_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg118_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
   MUX_Subtract2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract2_impl_0_LUT_out,
                 oMux => MUX_Subtract2_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_0_out,
                 Y => Delay1No146_out);

Delay3No_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast <= Delay3No_out;
SharedReg58_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg58_out;
   MUX_Subtract2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract2_impl_1_LUT_out,
                 oMux => MUX_Subtract2_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Subtract3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_impl_out,
                 X => Delay1No148_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast);

Delay3No5_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast <= Delay3No5_out;
Delay47No_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast <= Delay47No_out;
   MUX_Subtract3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No5_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay47No_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract3_impl_0_LUT_out,
                 oMux => MUX_Subtract3_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_0_out,
                 Y => Delay1No148_out);

Delay2No16_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast <= Delay2No16_out;
SharedReg149_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg149_out;
   MUX_Subtract3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No16_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract3_impl_1_LUT_out,
                 oMux => MUX_Subtract3_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Add112_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Add112_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Add112_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add112_impl_out,
                 X => Delay1No150_out_to_Add112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Add112_impl_parent_implementedSystem_port_1_cast);

Delay13No_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast <= Delay13No_out;
Delay79No1_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast <= Delay79No1_out;
   MUX_Add112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay13No_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay79No1_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add112_impl_0_LUT_out,
                 oMux => MUX_Add112_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_0_out,
                 Y => Delay1No150_out);

SharedReg62_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg144_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg144_out;
   MUX_Add112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg144_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add112_impl_1_LUT_out,
                 oMux => MUX_Add112_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Add12_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Add12_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Add12_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_impl_out,
                 X => Delay1No152_out_to_Add12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Add12_impl_parent_implementedSystem_port_1_cast);

Delay63No_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast <= Delay63No_out;
SharedReg169_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast <= SharedReg169_out;
   MUX_Add12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay63No_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg169_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add12_impl_0_LUT_out,
                 oMux => MUX_Add12_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_impl_0_out,
                 Y => Delay1No152_out);

SharedReg143_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg64_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg64_out;
   MUX_Add12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg64_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add12_impl_1_LUT_out,
                 oMux => MUX_Add12_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Add15_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Add15_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Add15_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_impl_out,
                 X => Delay1No154_out_to_Add15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Add15_impl_parent_implementedSystem_port_1_cast);

Delay81No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast <= Delay81No_out;
Delay33No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast <= Delay33No_out;
   MUX_Add15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay81No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay33No_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add15_impl_0_LUT_out,
                 oMux => MUX_Add15_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_0_out,
                 Y => Delay1No154_out);

SharedReg66_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg146_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Add15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add15_impl_1_LUT_out,
                 oMux => MUX_Add15_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Add4_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Add4_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Add4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add4_impl_out,
                 X => Delay1No156_out_to_Add4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Add4_impl_parent_implementedSystem_port_1_cast);

Delay5No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast <= Delay5No_out;
Delay30No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast <= Delay30No_out;
   MUX_Add4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay30No_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add4_impl_0_LUT_out,
                 oMux => MUX_Add4_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add4_impl_0_out,
                 Y => Delay1No156_out);

SharedReg68_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg170_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg170_out;
   MUX_Add4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add4_impl_1_LUT_out,
                 oMux => MUX_Add4_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add4_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Add7_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Add7_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Add7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_impl_out,
                 X => Delay1No158_out_to_Add7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Add7_impl_parent_implementedSystem_port_1_cast);

Delay5No8_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast <= Delay5No8_out;
Delay35No_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast <= Delay35No_out;
   MUX_Add7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No8_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay35No_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add7_impl_0_LUT_out,
                 oMux => MUX_Add7_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_0_out,
                 Y => Delay1No158_out);

SharedReg70_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg171_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg171_out;
   MUX_Add7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add7_impl_1_LUT_out,
                 oMux => MUX_Add7_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Add9_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Add9_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Add9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_impl_out,
                 X => Delay1No160_out_to_Add9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Add9_impl_parent_implementedSystem_port_1_cast);

Delay5No15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast <= Delay5No15_out;
Delay51No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast <= Delay51No_out;
   MUX_Add9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No15_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay51No_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add9_impl_0_LUT_out,
                 oMux => MUX_Add9_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_0_out,
                 Y => Delay1No160_out);

SharedReg72_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg172_out;
   MUX_Add9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add9_impl_1_LUT_out,
                 oMux => MUX_Add9_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_1_out,
                 Y => Delay1No161_out);
   Constant1_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_impl_out);

Delay1No162_out_to_Divide_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Divide_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Divide_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_impl_out,
                 X => Delay1No162_out_to_Divide_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Divide_impl_parent_implementedSystem_port_1_cast);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay107No1_out,
                 Y => Delay1No162_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product116_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product116_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product116_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product116_impl_out,
                 X => Delay1No164_out_to_Product116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product116_impl_parent_implementedSystem_port_1_cast);

SharedReg26_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg134_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg134_out;
   MUX_Product116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product116_impl_0_LUT_out,
                 oMux => MUX_Product116_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_0_out,
                 Y => Delay1No164_out);

SharedReg15_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg182_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product116_impl_1_LUT_out,
                 oMux => MUX_Product116_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product10_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product10_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product10_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_impl_out,
                 X => Delay1No166_out_to_Product10_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product10_impl_parent_implementedSystem_port_1_cast);

Delay2No43_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast <= Delay2No43_out;
SharedReg146_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product10_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No43_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product10_impl_0_LUT_out,
                 oMux => MUX_Product10_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_0_out,
                 Y => Delay1No166_out);

SharedReg149_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg185_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast <= SharedReg185_out;
   MUX_Product10_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product10_impl_1_LUT_out,
                 oMux => MUX_Product10_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product13_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product13_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product13_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_impl_out,
                 X => Delay1No168_out_to_Product13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product13_impl_parent_implementedSystem_port_1_cast);

SharedReg135_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg135_out;
Delay2No39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast <= Delay2No39_out;
   MUX_Product13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay2No39_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product13_impl_0_LUT_out,
                 oMux => MUX_Product13_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_0_out,
                 Y => Delay1No168_out);

SharedReg182_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg187_out;
   MUX_Product13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product13_impl_1_LUT_out,
                 oMux => MUX_Product13_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product16_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product16_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product16_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product16_impl_out,
                 X => Delay1No170_out_to_Product16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product16_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg146_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product16_impl_0_LUT_out,
                 oMux => MUX_Product16_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_0_out,
                 Y => Delay1No170_out);

SharedReg30_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg175_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Product16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product16_impl_1_LUT_out,
                 oMux => MUX_Product16_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product18_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product18_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product18_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_impl_out,
                 X => Delay1No172_out_to_Product18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product18_impl_parent_implementedSystem_port_1_cast);

Delay3No15_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast <= Delay3No15_out;
SharedReg151_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg151_out;
   MUX_Product18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No15_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product18_impl_0_LUT_out,
                 oMux => MUX_Product18_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_impl_0_out,
                 Y => Delay1No172_out);

SharedReg14_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg180_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg180_out;
   MUX_Product18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg180_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product18_impl_1_LUT_out,
                 oMux => MUX_Product18_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product19_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product19_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product19_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_impl_out,
                 X => Delay1No174_out_to_Product19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product19_impl_parent_implementedSystem_port_1_cast);

SharedReg159_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast <= SharedReg159_out;
SharedReg146_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product19_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg159_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product19_impl_0_LUT_out,
                 oMux => MUX_Product19_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_impl_0_out,
                 Y => Delay1No174_out);

SharedReg151_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg182_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product19_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product19_impl_1_LUT_out,
                 oMux => MUX_Product19_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product21_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product21_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product21_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_impl_out,
                 X => Delay1No176_out_to_Product21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product21_impl_parent_implementedSystem_port_1_cast);

SharedReg25_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg133_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast <= SharedReg133_out;
   MUX_Product21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg133_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product21_impl_0_LUT_out,
                 oMux => MUX_Product21_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_0_out,
                 Y => Delay1No176_out);

SharedReg149_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg175_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Product21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product21_impl_1_LUT_out,
                 oMux => MUX_Product21_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product23_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product23_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product23_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_impl_out,
                 X => Delay1No178_out_to_Product23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product23_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg103_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast <= SharedReg103_out;
   MUX_Product23_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg103_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product23_impl_0_LUT_out,
                 oMux => MUX_Product23_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_0_out,
                 Y => Delay1No178_out);

SharedReg15_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg188_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast <= SharedReg188_out;
   MUX_Product23_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product23_impl_1_LUT_out,
                 oMux => MUX_Product23_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product28_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product28_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product28_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_impl_out,
                 X => Delay1No180_out_to_Product28_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product28_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg156_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
   MUX_Product28_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product28_impl_0_LUT_out,
                 oMux => MUX_Product28_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_impl_0_out,
                 Y => Delay1No180_out);

SharedReg10_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg182_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product28_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product28_impl_1_LUT_out,
                 oMux => MUX_Product28_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product31_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product31_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product31_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_impl_out,
                 X => Delay1No182_out_to_Product31_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product31_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg160_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast <= SharedReg160_out;
   MUX_Product31_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg160_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product31_impl_0_LUT_out,
                 oMux => MUX_Product31_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_0_out,
                 Y => Delay1No182_out);

SharedReg26_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg182_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product31_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product31_impl_1_LUT_out,
                 oMux => MUX_Product31_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product34_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product34_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product34_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product34_impl_out,
                 X => Delay1No184_out_to_Product34_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product34_impl_parent_implementedSystem_port_1_cast);

SharedReg26_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg162_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_2_cast <= SharedReg162_out;
   MUX_Product34_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg162_out_to_MUX_Product34_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product34_impl_0_LUT_out,
                 oMux => MUX_Product34_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_impl_0_out,
                 Y => Delay1No184_out);

SharedReg10_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg175_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Product34_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product34_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product34_impl_1_LUT_out,
                 oMux => MUX_Product34_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product34_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product4_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product4_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_impl_out,
                 X => Delay1No186_out_to_Product4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product4_impl_parent_implementedSystem_port_1_cast);

SharedReg158_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg158_out;
SharedReg151_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg151_out;
   MUX_Product4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg158_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product4_impl_0_LUT_out,
                 oMux => MUX_Product4_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_0_out,
                 Y => Delay1No186_out);

SharedReg149_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg182_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Product4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product4_impl_1_LUT_out,
                 oMux => MUX_Product4_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product40_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product40_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product40_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product40_impl_out,
                 X => Delay1No188_out_to_Product40_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product40_impl_parent_implementedSystem_port_1_cast);

SharedReg21_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg163_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast <= SharedReg163_out;
   MUX_Product40_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg163_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product40_impl_0_LUT_out,
                 oMux => MUX_Product40_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product40_impl_0_out,
                 Y => Delay1No188_out);

SharedReg175_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg15_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product40_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product40_impl_1_LUT_out,
                 oMux => MUX_Product40_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product40_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product43_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product43_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product43_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product43_impl_out,
                 X => Delay1No190_out_to_Product43_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product43_impl_parent_implementedSystem_port_1_cast);

SharedReg164_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg121_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
   MUX_Product43_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product43_impl_0_LUT_out,
                 oMux => MUX_Product43_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product43_impl_0_out,
                 Y => Delay1No190_out);

SharedReg175_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg184_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast <= SharedReg184_out;
   MUX_Product43_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product43_impl_1_LUT_out,
                 oMux => MUX_Product43_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product43_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product44_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product44_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product44_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product44_impl_out,
                 X => Delay1No192_out_to_Product44_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product44_impl_parent_implementedSystem_port_1_cast);

SharedReg168_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast <= SharedReg168_out;
SharedReg122_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
   MUX_Product44_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product44_impl_0_LUT_out,
                 oMux => MUX_Product44_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product44_impl_0_out,
                 Y => Delay1No192_out);

SharedReg180_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast <= SharedReg180_out;
SharedReg179_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast <= SharedReg179_out;
   MUX_Product44_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg180_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product44_impl_1_LUT_out,
                 oMux => MUX_Product44_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product44_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product47_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product47_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product47_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product47_impl_out,
                 X => Delay1No194_out_to_Product47_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product47_impl_parent_implementedSystem_port_1_cast);

Delay1No226_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_1_cast <= Delay1No226_out;
SharedReg116_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_2_cast <= SharedReg116_out;
   MUX_Product47_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay1No226_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Product47_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product47_impl_0_LUT_out,
                 oMux => MUX_Product47_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product47_impl_0_out,
                 Y => Delay1No194_out);

SharedReg180_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_1_cast <= SharedReg180_out;
SharedReg173_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
   MUX_Product47_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg180_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product47_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product47_impl_1_LUT_out,
                 oMux => MUX_Product47_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product47_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product49_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product49_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product49_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product49_impl_out,
                 X => Delay1No196_out_to_Product49_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product49_impl_parent_implementedSystem_port_1_cast);

Delay1No227_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast <= Delay1No227_out;
SharedReg166_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast <= SharedReg166_out;
   MUX_Product49_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay1No227_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product49_impl_0_LUT_out,
                 oMux => MUX_Product49_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product49_impl_0_out,
                 Y => Delay1No196_out);

SharedReg182_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg173_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
   MUX_Product49_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product49_impl_1_LUT_out,
                 oMux => MUX_Product49_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product49_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product6_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product6_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_impl_out,
                 X => Delay1No198_out_to_Product6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product6_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
Delay1No228_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast <= Delay1No228_out;
   MUX_Product6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No228_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product6_impl_0_LUT_out,
                 oMux => MUX_Product6_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_0_out,
                 Y => Delay1No198_out);

SharedReg11_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg173_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg173_out;
   MUX_Product6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product6_impl_1_LUT_out,
                 oMux => MUX_Product6_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_1_out,
                 Y => Delay1No199_out);
   Constant_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_impl_out);

   Delay5No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_out,
                 Y => Delay5No_out);

   Delay12No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => Delay12No_out);

   Delay11No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => Delay11No_out);

   Delay5No8_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_out,
                 Y => Delay5No8_out);

   Delay12No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => Delay12No1_out);

   Delay11No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => Delay11No1_out);

   Delay11No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => Delay11No2_out);

   Delay5No15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_out,
                 Y => Delay5No15_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_out,
                 Y => Delay1No226_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_out,
                 Y => Delay1No227_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_out,
                 Y => Delay1No228_out);

   Delay90No_instance: Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=88 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => Delay90No_out);

   Delay93No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay93No_out);

   Delay93No1_instance: Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=90 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => Delay93No1_out);

   Delay3No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay3No_out);

   Delay79No_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => Delay79No_out);

   Delay97No_instance: Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=95 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => Delay97No_out);

   Delay97No1_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => Delay97No1_out);

   Delay2No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay2No16_out);

   Delay94No_instance: Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=93 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => Delay94No_out);

   Delay2No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => Delay2No17_out);

   Delay89No_instance: Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=87 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay89No_out);

   Delay18No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => Delay18No_out);

   Delay23No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay23No_out);

   Delay9No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => Delay9No_out);

   Delay6No10_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay6No10_out);

   Delay12No2_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay12No2_out);

   Delay7No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay7No2_out);

   Delay15No_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => Delay15No_out);

   Delay3No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => Delay3No5_out);

   Delay12No3_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => Delay12No3_out);

   Delay8No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => Delay8No1_out);

   Delay20No_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => Delay20No_out);

   Delay7No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => Delay7No4_out);

   Delay10No7_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => Delay10No7_out);

   Delay8No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay8No2_out);

   Delay3No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => Delay3No7_out);

   Delay6No12_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => Delay6No12_out);

   Delay8No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => Delay8No3_out);

   Delay103No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => Delay103No_out);

   Delay107No_instance: Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=105 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay107No_out);

   Delay89No1_instance: Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=82 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => Delay89No1_out);

   Delay89No2_instance: Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=82 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => Delay89No2_out);

   Delay18No1_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay18No1_out);

   Delay22No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => Delay22No_out);

   Delay14No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => Delay14No_out);

   Delay3No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay3No11_out);

   Delay11No3_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => Delay11No3_out);

   Delay15No2_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => Delay15No2_out);

   Delay12No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => Delay12No4_out);

   Delay17No_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => Delay17No_out);

   Delay2No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => Delay2No35_out);

   Delay3No13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => Delay3No13_out);

   Delay96No_instance: Delay_34_DelayLength_93_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=93 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => Delay96No_out);

   Delay107No1_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_impl_out,
                 Y => Delay107No1_out);

   Delay63No_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay63No_out);

   Delay61No_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => Delay61No_out);

   Delay65No_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => Delay65No_out);

   Delay81No_instance: Delay_34_DelayLength_71_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=71 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => Delay81No_out);

   Delay51No_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => Delay51No_out);

   Delay2No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => Delay2No36_out);

   Delay44No_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => Delay44No_out);

   Delay2No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => Delay2No38_out);

   Delay47No_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => Delay47No_out);

   Delay2No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => Delay2No39_out);

   Delay35No_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => Delay35No_out);

   Delay31No_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => Delay31No_out);

   Delay3No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay3No15_out);

   Delay33No_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => Delay33No_out);

   Delay30No_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => Delay30No_out);

   Delay25No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => Delay25No1_out);

   Delay13No_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => Delay13No_out);

   Delay2No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => Delay2No42_out);

   Delay79No1_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => Delay79No1_out);

   Delay2No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => Delay2No43_out);

   Delay21No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => Delay21No_out);

   MUX_Add24_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add24_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add24_impl_0_LUT_out);

   MUX_Add24_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add24_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add24_impl_1_LUT_out);

   MUX_Add61_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add61_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add61_impl_0_LUT_out);

   MUX_Add61_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add61_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add61_impl_1_LUT_out);

   MUX_Product74_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product74_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product74_impl_0_LUT_out);

   MUX_Product74_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product74_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product74_impl_1_LUT_out);

   MUX_Product76_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product76_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product76_impl_0_LUT_out);

   MUX_Product76_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product76_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product76_impl_1_LUT_out);

   MUX_Product77_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product77_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product77_impl_0_LUT_out);

   MUX_Product77_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product77_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product77_impl_1_LUT_out);

   MUX_Product81_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product81_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product81_impl_0_LUT_out);

   MUX_Product81_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product81_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product81_impl_1_LUT_out);

   MUX_Product84_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product84_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product84_impl_0_LUT_out);

   MUX_Product84_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product84_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product84_impl_1_LUT_out);

   MUX_Product86_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product86_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product86_impl_0_LUT_out);

   MUX_Product86_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product86_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product86_impl_1_LUT_out);

   MUX_Product87_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product87_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product87_impl_0_LUT_out);

   MUX_Product87_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product87_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product87_impl_1_LUT_out);

   MUX_Product88_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product88_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product88_impl_0_LUT_out);

   MUX_Product88_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product88_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product88_impl_1_LUT_out);

   MUX_Product94_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product94_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product94_impl_0_LUT_out);

   MUX_Product94_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product94_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product94_impl_1_LUT_out);

   MUX_Product97_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product97_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product97_impl_0_LUT_out);

   MUX_Product97_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product97_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product97_impl_1_LUT_out);

   MUX_Product98_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product98_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product98_impl_0_LUT_out);

   MUX_Product98_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product98_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product98_impl_1_LUT_out);

   MUX_Product99_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product99_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product99_impl_0_LUT_out);

   MUX_Product99_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product99_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product99_impl_1_LUT_out);

   MUX_Subtract2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract2_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Subtract2_impl_0_LUT_out);

   MUX_Subtract2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract2_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Subtract2_impl_1_LUT_out);

   MUX_Subtract3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract3_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Subtract3_impl_0_LUT_out);

   MUX_Subtract3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract3_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Subtract3_impl_1_LUT_out);

   MUX_Add112_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add112_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add112_impl_0_LUT_out);

   MUX_Add112_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add112_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add112_impl_1_LUT_out);

   MUX_Add12_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add12_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add12_impl_0_LUT_out);

   MUX_Add12_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add12_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add12_impl_1_LUT_out);

   MUX_Add15_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add15_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add15_impl_0_LUT_out);

   MUX_Add15_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add15_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add15_impl_1_LUT_out);

   MUX_Add4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add4_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add4_impl_0_LUT_out);

   MUX_Add4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add4_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add4_impl_1_LUT_out);

   MUX_Add7_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add7_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add7_impl_0_LUT_out);

   MUX_Add7_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add7_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add7_impl_1_LUT_out);

   MUX_Add9_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add9_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add9_impl_0_LUT_out);

   MUX_Add9_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add9_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Add9_impl_1_LUT_out);

   MUX_Product116_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product116_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product116_impl_0_LUT_out);

   MUX_Product116_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product116_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product116_impl_1_LUT_out);

   MUX_Product10_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product10_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product10_impl_0_LUT_out);

   MUX_Product10_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product10_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product10_impl_1_LUT_out);

   MUX_Product13_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product13_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product13_impl_0_LUT_out);

   MUX_Product13_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product13_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product13_impl_1_LUT_out);

   MUX_Product16_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product16_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product16_impl_0_LUT_out);

   MUX_Product16_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product16_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product16_impl_1_LUT_out);

   MUX_Product18_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product18_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product18_impl_0_LUT_out);

   MUX_Product18_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product18_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product18_impl_1_LUT_out);

   MUX_Product19_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product19_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product19_impl_0_LUT_out);

   MUX_Product19_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product19_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product19_impl_1_LUT_out);

   MUX_Product21_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product21_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product21_impl_0_LUT_out);

   MUX_Product21_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product21_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product21_impl_1_LUT_out);

   MUX_Product23_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product23_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product23_impl_0_LUT_out);

   MUX_Product23_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product23_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product23_impl_1_LUT_out);

   MUX_Product28_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product28_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product28_impl_0_LUT_out);

   MUX_Product28_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product28_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product28_impl_1_LUT_out);

   MUX_Product31_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product31_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product31_impl_0_LUT_out);

   MUX_Product31_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product31_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product31_impl_1_LUT_out);

   MUX_Product34_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product34_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product34_impl_0_LUT_out);

   MUX_Product34_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product34_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product34_impl_1_LUT_out);

   MUX_Product4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product4_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product4_impl_0_LUT_out);

   MUX_Product4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product4_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product4_impl_1_LUT_out);

   MUX_Product40_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product40_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product40_impl_0_LUT_out);

   MUX_Product40_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product40_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product40_impl_1_LUT_out);

   MUX_Product43_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product43_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product43_impl_0_LUT_out);

   MUX_Product43_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product43_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product43_impl_1_LUT_out);

   MUX_Product44_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product44_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product44_impl_0_LUT_out);

   MUX_Product44_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product44_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product44_impl_1_LUT_out);

   MUX_Product47_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product47_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product47_impl_0_LUT_out);

   MUX_Product47_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product47_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product47_impl_1_LUT_out);

   MUX_Product49_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product49_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product49_impl_0_LUT_out);

   MUX_Product49_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product49_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product49_impl_1_LUT_out);

   MUX_Product6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product6_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product6_impl_0_LUT_out);

   MUX_Product6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product6_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount31_out,
                 Output => MUX_Product6_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_impl_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_impl_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_impl_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_impl_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_impl_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_impl_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_impl_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_impl_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_impl_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_impl_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_impl_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_impl_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_impl_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add19_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add20_impl_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add21_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=74 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add22_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_impl_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add61_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product1010_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product101_impl_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_impl_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product121_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product141_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product161_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product171_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product181_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product191_impl_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product241_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product271_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_impl_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product331_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product351_impl_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product411_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product412_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product57_impl_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product58_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product59_impl_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product60_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product64_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product65_impl_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product66_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product72_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product74_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product76_impl_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product77_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product81_impl_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product84_impl_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product86_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product87_impl_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product88_impl_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product94_impl_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product97_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product98_impl_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product99_impl_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract1_impl_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract11_impl_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_impl_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add112_impl_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_impl_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add4_impl_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_impl_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_impl_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_impl_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product116_impl_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_impl_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product16_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_impl_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_impl_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_impl_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_impl_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product34_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_impl_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product40_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product43_impl_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product44_impl_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product47_impl_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product49_impl_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_impl_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_impl_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);
end architecture;

