--------------------------------------------------------------------------------
--                         ModuloCounter_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_2_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of ModuloCounter_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(0 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 1 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2292563
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2292563 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2292563 is
signal XX_m2292564 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2292564 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2292564 <= X ;
   YY_m2292564 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2292567
--                   (IntAdderClassical_33_f500_uid2292569)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2292567 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2292567 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2292563 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2292567 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2292563  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2292567  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2292874_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2292876)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2292874_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2292874_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2292879
--                  (IntAdderAlternative_27_f250_uid2292883)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2292879 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2292879 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2292886
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2292886 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2292886 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2292889
--                   (IntAdderClassical_34_f250_uid2292891)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2292889 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2292889 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2292874
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2292874 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2292874 is
   component FPAdd_8_23_uid2292874_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2292879 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2292886 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2292889 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2292874_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2292879  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2292886  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2292889  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2292874 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2292874  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2294641_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2294643)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2294641_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2294641_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2294646
--                  (IntAdderAlternative_27_f250_uid2294650)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2294646 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2294646 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2294653
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2294653 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2294653 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2294656
--                   (IntAdderClassical_34_f250_uid2294658)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2294656 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2294656 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2294641
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2294641 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2294641 is
   component FPAdd_8_23_uid2294641_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2294646 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2294653 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2294656 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2294641_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2294646  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2294653  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2294656  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2294641 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2294641  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 91 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      Y <= s90;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 92 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      Y <= s91;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 96 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      Y <= s95;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 74 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      Y <= s73;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 81 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      Y <= s80;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 82 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      Y <= s81;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 95 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      Y <= s94;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 90 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      Y <= s89;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 107 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      Y <= s106;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 64 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      Y <= s63;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 51 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      Y <= s50;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 76 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      Y <= s75;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 79 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      Y <= s78;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1 : in std_logic_vector(31 downto 0);
          R_U : in std_logic_vector(31 downto 0);
          R_V : in std_logic_vector(31 downto 0);
          R_W : in std_logic_vector(31 downto 0);
          Inv_11 : out std_logic_vector(31 downto 0);
          Inv_12 : out std_logic_vector(31 downto 0);
          Inv_13 : out std_logic_vector(31 downto 0);
          Inv_21 : out std_logic_vector(31 downto 0);
          Inv_22 : out std_logic_vector(31 downto 0);
          Inv_23 : out std_logic_vector(31 downto 0);
          Inv_31 : out std_logic_vector(31 downto 0);
          Inv_32 : out std_logic_vector(31 downto 0);
          Inv_33 : out std_logic_vector(31 downto 0);
          Inv_41 : out std_logic_vector(31 downto 0);
          Inv_42 : out std_logic_vector(31 downto 0);
          Inv_43 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_2_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(0 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount21_out : std_logic_vector(0 downto 0) := (others => '0');
signal Ldiff_UU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add151_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add210_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add27_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add27_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add29_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add29_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add29_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add31_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add31_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add51_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add51_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add51_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add61_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add71_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add71_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add71_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add81_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product101_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product101_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product101_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product121_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product121_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product141_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product141_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product151_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product151_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product151_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product171_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product171_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product171_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product181_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product181_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product212_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product212_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product212_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product241_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product251_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product251_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product251_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product261_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product261_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product261_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product271_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product271_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product271_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product361_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product361_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product361_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product401_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product401_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product401_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product412_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product412_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product412_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product431_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product431_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product471_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product471_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product471_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product481_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product491_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product491_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product512_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product512_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product59_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product61_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product63_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product65_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product65_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product65_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product66_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product67_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product72_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product73_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product73_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product73_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product76_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product77_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product77_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product77_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product81_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product81_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product81_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product82_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product82_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product82_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product83_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product83_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product83_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product84_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product84_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product84_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product87_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product87_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product87_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product90_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product90_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product90_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product91_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product91_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product91_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product93_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product93_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product93_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product96_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product96_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product96_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product98_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product98_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product98_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product99_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product99_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product99_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add211_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product115_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product115_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product29_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay66No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay81No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay46No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay49No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No448_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No449_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay31No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay29No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No454_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No456_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No457_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No458_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No459_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No460_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No461_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No464_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No16_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay82No_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay83No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No31_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No4_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay92No2_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add101_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add101_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No3_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add131_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add131_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add141_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add141_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add151_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add151_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No1_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No2_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add210_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add210_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No38_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay66No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No1_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay34No_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add29_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add29_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add31_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add31_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay46No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add51_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add51_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No34_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add61_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add61_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No24_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add71_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add71_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No2_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add81_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add81_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product113_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product113_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product101_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product101_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No17_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product121_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product121_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product141_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product141_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product151_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product151_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product171_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product171_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No22_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product181_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product181_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product212_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product212_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product221_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product221_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product241_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product241_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product251_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product251_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No18_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product261_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product261_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product271_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product271_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product312_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product312_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product321_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product321_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No13_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product361_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product361_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product401_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product401_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product412_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product412_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product431_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product431_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No20_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product471_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product471_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product481_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product481_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product491_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product491_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product512_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product512_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product54_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product54_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product55_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product55_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product59_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product59_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No22_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product61_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product61_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product63_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product63_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product65_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product65_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product66_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product66_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No23_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product67_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product67_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No15_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Product68_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Product68_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No16_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product72_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product72_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product73_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product73_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product76_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product76_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product77_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product77_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product81_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product81_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No29_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product82_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product82_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product83_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product83_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product84_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product84_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product87_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product87_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product90_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product90_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product91_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product91_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product93_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product93_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product96_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product96_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product98_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product98_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product99_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product99_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No11_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No18_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No15_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No23_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No4_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Subtract5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Subtract5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No12_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Add32_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Add32_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Add11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Add11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Add13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Add13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Add15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Add15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Add211_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Add211_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Add4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Add4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Add6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Add6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Add9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Add9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Divide_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Divide_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product115_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product115_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product10_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product10_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product14_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product14_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Product17_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Product17_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Product18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Product18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product213_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product213_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Product22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Product22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Product23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Product23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product26_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product26_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product28_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product28_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product29_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product29_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Product3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Product3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Product30_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Product30_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product31_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product31_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product32_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product32_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product33_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product33_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product34_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product34_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Product36_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Product36_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Product37_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Product37_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product38_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product38_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Product43_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Product43_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Product44_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Product44_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Product45_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Product45_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Product46_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Product46_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product47_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product47_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product48_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product48_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Product49_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Product49_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Product5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Product5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Product50_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Product50_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Product7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Product7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Subtract_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Subtract_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount21_instance: ModuloCounter_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount21_out);
Ldiff_UU_del_1_IEEE <= Ldiff_UU_del_1;
   Ldiff_UU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_out,
                 X => Ldiff_UU_del_1_IEEE);
Ldiff_UV_del_1_IEEE <= Ldiff_UV_del_1;
   Ldiff_UV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_out,
                 X => Ldiff_UV_del_1_IEEE);
Ldiff_UW_del_1_IEEE <= Ldiff_UW_del_1;
   Ldiff_UW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_out,
                 X => Ldiff_UW_del_1_IEEE);
Ldiff_VU_del_1_IEEE <= Ldiff_VU_del_1;
   Ldiff_VU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_out,
                 X => Ldiff_VU_del_1_IEEE);
Ldiff_VV_del_1_IEEE <= Ldiff_VV_del_1;
   Ldiff_VV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_out,
                 X => Ldiff_VV_del_1_IEEE);
Ldiff_VW_del_1_IEEE <= Ldiff_VW_del_1;
   Ldiff_VW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_out,
                 X => Ldiff_VW_del_1_IEEE);
Ldiff_WU_del_1_IEEE <= Ldiff_WU_del_1;
   Ldiff_WU_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_out,
                 X => Ldiff_WU_del_1_IEEE);
Ldiff_WV_del_1_IEEE <= Ldiff_WV_del_1;
   Ldiff_WV_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_out,
                 X => Ldiff_WV_del_1_IEEE);
Ldiff_WW_del_1_IEEE <= Ldiff_WW_del_1;
   Ldiff_WW_del_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_out,
                 X => Ldiff_WW_del_1_IEEE);
R_U_IEEE <= R_U;
   R_U_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_out,
                 X => R_U_IEEE);
R_V_IEEE <= R_V;
   R_V_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_out,
                 X => R_V_IEEE);
R_W_IEEE <= R_W;
   R_W_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_out,
                 X => R_W_IEEE);

Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_impl_out,
                 X => Delay1No_out_to_Product108_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_impl_parent_implementedSystem_port_1_cast);

Delay5No16_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast <= Delay5No16_out;
SharedReg117_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product108_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No16_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product108_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product108_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_impl_0_out,
                 Y => Delay1No_out);

SharedReg61_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
Delay92No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast <= Delay92No_out;
   MUX_Product108_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay92No_out_to_MUX_Product108_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product108_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product110_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_impl_out,
                 X => Delay1No2_out_to_Product110_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product110_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg117_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product110_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product110_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product110_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_impl_0_out,
                 Y => Delay1No2_out);

SharedReg131_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
Delay97No2_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast <= Delay97No2_out;
   MUX_Product110_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No2_out_to_MUX_Product110_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product110_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product109_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_impl_out,
                 X => Delay1No4_out_to_Product109_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product109_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg117_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product109_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product109_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product109_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_impl_0_out,
                 Y => Delay1No4_out);

SharedReg16_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
Delay82No_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast <= Delay82No_out;
   MUX_Product109_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay82No_out_to_MUX_Product109_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product109_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product111_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_impl_out,
                 X => Delay1No6_out_to_Product111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product111_impl_parent_implementedSystem_port_1_cast);

SharedReg109_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast <= SharedReg109_out;
SharedReg117_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg109_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product111_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_0_out,
                 Y => Delay1No6_out);

SharedReg136_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
Delay83No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast <= Delay83No_out;
   MUX_Product111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay83No_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product111_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product210_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_impl_out,
                 X => Delay1No8_out_to_Product210_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product210_impl_parent_implementedSystem_port_1_cast);

Delay2No31_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast <= Delay2No31_out;
SharedReg117_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product210_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No31_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product210_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_0_out,
                 Y => Delay1No8_out);

SharedReg133_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
Delay97No3_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast <= Delay97No3_out;
   MUX_Product210_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No3_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product210_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product310_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_impl_out,
                 X => Delay1No10_out_to_Product310_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product310_impl_parent_implementedSystem_port_1_cast);

SharedReg110_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg117_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product310_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product310_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_0_out,
                 Y => Delay1No10_out);

SharedReg136_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
Delay97No4_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast <= Delay97No4_out;
   MUX_Product310_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No4_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product310_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product410_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_impl_out,
                 X => Delay1No12_out_to_Product410_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product410_impl_parent_implementedSystem_port_1_cast);

SharedReg111_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg117_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product410_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product410_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product410_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_impl_0_out,
                 Y => Delay1No12_out);

SharedReg136_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
Delay92No2_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast <= Delay92No2_out;
   MUX_Product410_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay92No2_out_to_MUX_Product410_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product410_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product510_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_impl_out,
                 X => Delay1No14_out_to_Product510_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product510_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg117_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product510_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product510_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product510_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_impl_0_out,
                 Y => Delay1No14_out);

SharedReg133_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
Delay95No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast <= Delay95No_out;
   MUX_Product510_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay95No_out_to_MUX_Product510_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product510_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product610_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_impl_out,
                 X => Delay1No16_out_to_Product610_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product610_impl_parent_implementedSystem_port_1_cast);

Delay2No17_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast <= Delay2No17_out;
SharedReg117_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product610_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No17_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product610_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product610_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_impl_0_out,
                 Y => Delay1No16_out);

SharedReg133_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
Delay97No_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast <= Delay97No_out;
   MUX_Product610_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No_out_to_MUX_Product610_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product610_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product710_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_impl_out,
                 X => Delay1No18_out_to_Product710_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product710_impl_parent_implementedSystem_port_1_cast);

Delay6No12_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast <= Delay6No12_out;
SharedReg117_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product710_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No12_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product710_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product710_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_impl_0_out,
                 Y => Delay1No18_out);

SharedReg61_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
Delay97No1_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast <= Delay97No1_out;
   MUX_Product710_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No1_out_to_MUX_Product710_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product710_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product810_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_impl_out,
                 X => Delay1No20_out_to_Product810_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product810_impl_parent_implementedSystem_port_1_cast);

SharedReg66_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg117_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product810_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product810_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product810_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_impl_0_out,
                 Y => Delay1No20_out);

SharedReg8_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg44_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast <= SharedReg44_out;
   MUX_Product810_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg44_out_to_MUX_Product810_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product810_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product910_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_impl_out,
                 X => Delay1No22_out_to_Product910_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product910_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg117_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Product910_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product910_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product910_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_impl_0_out,
                 Y => Delay1No22_out);

SharedReg131_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
Delay75No_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast <= Delay75No_out;
   MUX_Product910_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay75No_out_to_MUX_Product910_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product910_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_impl_1_out,
                 Y => Delay1No23_out);
   Inv_11_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_IEEE,
                 X => Delay1No24_out);
Inv_11 <= Inv_11_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => Delay1No24_out);
   Inv_12_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_IEEE,
                 X => Delay1No25_out);
Inv_12 <= Inv_12_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => Delay1No25_out);
   Inv_13_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_IEEE,
                 X => Delay1No26_out);
Inv_13 <= Inv_13_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => Delay1No26_out);
   Inv_21_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_IEEE,
                 X => Delay1No27_out);
Inv_21 <= Inv_21_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => Delay1No27_out);
   Inv_22_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_IEEE,
                 X => Delay1No28_out);
Inv_22 <= Inv_22_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => Delay1No28_out);
   Inv_23_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_IEEE,
                 X => Delay1No29_out);
Inv_23 <= Inv_23_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => Delay1No29_out);
   Inv_31_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_IEEE,
                 X => Delay1No30_out);
Inv_31 <= Inv_31_IEEE;

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay1No30_out);
   Inv_32_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_IEEE,
                 X => Delay1No31_out);
Inv_32 <= Inv_32_IEEE;

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => Delay1No31_out);
   Inv_33_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_IEEE,
                 X => Delay1No32_out);
Inv_33 <= Inv_33_IEEE;

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => Delay1No32_out);
   Inv_41_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_IEEE,
                 X => Delay1No33_out);
Inv_41 <= Inv_41_IEEE;

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => Delay1No33_out);
   Inv_42_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_IEEE,
                 X => Delay1No34_out);
Inv_42 <= Inv_42_IEEE;

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay1No34_out);
   Inv_43_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_IEEE,
                 X => Delay1No35_out);
Inv_43 <= Inv_43_IEEE;

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add30_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_impl_out,
                 X => Delay1No36_out_to_Add30_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add30_impl_parent_implementedSystem_port_1_cast);

SharedReg82_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast <= SharedReg82_out;
Delay17No_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast <= Delay17No_out;
   MUX_Add30_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg82_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay17No_out_to_MUX_Add30_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add30_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_impl_0_out,
                 Y => Delay1No36_out);

SharedReg94_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
   MUX_Add30_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Add30_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add30_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add101_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add101_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add101_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_impl_out,
                 X => Delay1No38_out_to_Add101_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add101_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg87_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast <= SharedReg87_out;
   MUX_Add101_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Add101_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add101_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_impl_0_out,
                 Y => Delay1No38_out);

SharedReg83_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg88_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast <= SharedReg88_out;
   MUX_Add101_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg88_out_to_MUX_Add101_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add101_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add111_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add111_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add111_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_impl_out,
                 X => Delay1No40_out_to_Add111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add111_impl_parent_implementedSystem_port_1_cast);

Delay9No_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast <= Delay9No_out;
Delay17No3_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast <= Delay17No3_out;
   MUX_Add111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay9No_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay17No3_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add111_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_0_out,
                 Y => Delay1No40_out);

SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg116_out;
SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg116_out;
   MUX_Add111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add111_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add131_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add131_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add131_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_impl_out,
                 X => Delay1No42_out_to_Add131_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add131_impl_parent_implementedSystem_port_1_cast);

Delay7No2_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast <= Delay7No2_out;
SharedReg107_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast <= SharedReg107_out;
   MUX_Add131_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No2_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg107_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add131_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_0_out,
                 Y => Delay1No42_out);

Delay2No36_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast <= Delay2No36_out;
SharedReg108_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
   MUX_Add131_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No36_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add131_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add141_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add141_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add141_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_impl_out,
                 X => Delay1No44_out_to_Add141_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add141_impl_parent_implementedSystem_port_1_cast);

SharedReg91_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_1_cast <= SharedReg91_out;
Delay18No_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_2_cast <= Delay18No_out;
   MUX_Add141_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay18No_out_to_MUX_Add141_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add141_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_impl_0_out,
                 Y => Delay1No44_out);

SharedReg92_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg55_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_2_cast <= SharedReg55_out;
   MUX_Add141_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Add141_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add141_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add151_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add151_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add151_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add151_impl_out,
                 X => Delay1No46_out_to_Add151_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add151_impl_parent_implementedSystem_port_1_cast);

Delay7No3_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_1_cast <= Delay7No3_out;
Delay4No_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_2_cast <= Delay4No_out;
   MUX_Add151_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No3_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No_out_to_MUX_Add151_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add151_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_impl_0_out,
                 Y => Delay1No46_out);

SharedReg115_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
Delay4No1_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_2_cast <= Delay4No1_out;
   MUX_Add151_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No1_out_to_MUX_Add151_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add151_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add16_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_impl_out,
                 X => Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
Delay20No_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast <= Delay20No_out;
   MUX_Add16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay20No_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add16_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_0_out,
                 Y => Delay1No48_out);

SharedReg96_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg113_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg113_out;
   MUX_Add16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg113_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add16_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add18_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add18_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add18_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_impl_out,
                 X => Delay1No50_out_to_Add18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add18_impl_parent_implementedSystem_port_1_cast);

SharedReg102_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg102_out;
SharedReg71_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg71_out;
   MUX_Add18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg102_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add18_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_0_out,
                 Y => Delay1No50_out);

Delay9No1_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast <= Delay9No1_out;
SharedReg72_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
   MUX_Add18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay9No1_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add18_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add19_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add19_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add19_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add19_impl_out,
                 X => Delay1No52_out_to_Add19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add19_impl_parent_implementedSystem_port_1_cast);

Delay15No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast <= Delay15No_out;
Delay17No2_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast <= Delay17No2_out;
   MUX_Add19_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay15No_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay17No2_out_to_MUX_Add19_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add19_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_impl_0_out,
                 Y => Delay1No52_out);

Delay2No11_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast <= Delay2No11_out;
SharedReg115_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast <= SharedReg115_out;
   MUX_Add19_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No11_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg115_out_to_MUX_Add19_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add19_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add210_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add210_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add210_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add210_impl_out,
                 X => Delay1No54_out_to_Add210_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add210_impl_parent_implementedSystem_port_1_cast);

SharedReg40_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
Delay14No_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_2_cast <= Delay14No_out;
   MUX_Add210_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay14No_out_to_MUX_Add210_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add210_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_impl_0_out,
                 Y => Delay1No54_out);

SharedReg68_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
Delay1No405_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_2_cast <= Delay1No405_out;
   MUX_Add210_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No405_out_to_MUX_Add210_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add210_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add20_impl_out,
                 X => Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast);

Delay19No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast <= Delay19No_out;
Delay64No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast <= Delay64No_out;
   MUX_Add20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay19No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay64No_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add20_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_0_out,
                 Y => Delay1No56_out);

Delay2No38_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast <= Delay2No38_out;
Delay1No420_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast <= Delay1No420_out;
   MUX_Add20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No38_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No420_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add20_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add21_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add21_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add21_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add21_impl_out,
                 X => Delay1No58_out_to_Add21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add21_impl_parent_implementedSystem_port_1_cast);

Delay25No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast <= Delay25No_out;
Delay66No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast <= Delay66No_out;
   MUX_Add21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay25No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay66No_out_to_MUX_Add21_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add21_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_impl_0_out,
                 Y => Delay1No58_out);

Delay2No13_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast <= Delay2No13_out;
Delay1No408_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast <= Delay1No408_out;
   MUX_Add21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No13_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No408_out_to_MUX_Add21_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add21_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add23_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add23_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add23_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_impl_out,
                 X => Delay1No60_out_to_Add23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add23_impl_parent_implementedSystem_port_1_cast);

SharedReg108_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_1_cast <= SharedReg108_out;
Delay76No_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_2_cast <= Delay76No_out;
   MUX_Add23_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg108_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay76No_out_to_MUX_Add23_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add23_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_impl_0_out,
                 Y => Delay1No60_out);

SharedReg45_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_1_cast <= SharedReg45_out;
Delay1No410_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_2_cast <= Delay1No410_out;
   MUX_Add23_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg45_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No410_out_to_MUX_Add23_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add23_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add24_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add24_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add24_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_impl_out,
                 X => Delay1No62_out_to_Add24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add24_impl_parent_implementedSystem_port_1_cast);

Delay11No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast <= Delay11No4_out;
Delay25No1_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast <= Delay25No1_out;
   MUX_Add24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No4_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay25No1_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add24_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_0_out,
                 Y => Delay1No62_out);

SharedReg112_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg112_out;
Delay1No413_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast <= Delay1No413_out;
   MUX_Add24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg112_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No413_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add24_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add27_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add27_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add27_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add27_impl_out,
                 X => Delay1No64_out_to_Add27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add27_impl_parent_implementedSystem_port_1_cast);

SharedReg36_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
Delay34No_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast <= Delay34No_out;
   MUX_Add27_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay34No_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add27_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add27_impl_0_out,
                 Y => Delay1No64_out);

SharedReg47_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast <= SharedReg47_out;
Delay1No415_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast <= Delay1No415_out;
   MUX_Add27_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No415_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add27_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add27_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add29_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add29_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add29_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add29_impl_out,
                 X => Delay1No66_out_to_Add29_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add29_impl_parent_implementedSystem_port_1_cast);

Delay17No1_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_1_cast <= Delay17No1_out;
Delay36No_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_2_cast <= Delay36No_out;
   MUX_Add29_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay17No1_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay36No_out_to_MUX_Add29_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add29_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add29_impl_0_out,
                 Y => Delay1No66_out);

SharedReg48_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
Delay1No417_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_2_cast <= Delay1No417_out;
   MUX_Add29_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No417_out_to_MUX_Add29_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add29_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add29_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add31_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add31_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add31_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add31_impl_out,
                 X => Delay1No68_out_to_Add31_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add31_impl_parent_implementedSystem_port_1_cast);

Delay12No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_1_cast <= Delay12No_out;
Delay46No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_2_cast <= Delay46No_out;
   MUX_Add31_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay46No_out_to_MUX_Add31_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add31_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add31_impl_0_out,
                 Y => Delay1No68_out);

SharedReg113_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_1_cast <= SharedReg113_out;
Delay1No466_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_2_cast <= Delay1No466_out;
   MUX_Add31_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No466_out_to_MUX_Add31_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add31_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add31_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add51_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add51_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add51_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add51_impl_out,
                 X => Delay1No70_out_to_Add51_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add51_impl_parent_implementedSystem_port_1_cast);

Delay11No1_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_1_cast <= Delay11No1_out;
Delay5No_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_2_cast <= Delay5No_out;
   MUX_Add51_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No1_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay5No_out_to_MUX_Add51_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add51_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add51_impl_0_out,
                 Y => Delay1No70_out);

Delay2No34_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_1_cast <= Delay2No34_out;
SharedReg124_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_2_cast <= SharedReg124_out;
   MUX_Add51_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No34_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Add51_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add51_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add51_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add61_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add61_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add61_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add61_impl_out,
                 X => Delay1No72_out_to_Add61_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add61_impl_parent_implementedSystem_port_1_cast);

SharedReg69_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast <= SharedReg69_out;
Delay5No7_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast <= Delay5No7_out;
   MUX_Add61_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay5No7_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add61_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_0_out,
                 Y => Delay1No72_out);

Delay2No24_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast <= Delay2No24_out;
SharedReg125_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast <= SharedReg125_out;
   MUX_Add61_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No24_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg125_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add61_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add71_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add71_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add71_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add71_impl_out,
                 X => Delay1No74_out_to_Add71_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add71_impl_parent_implementedSystem_port_1_cast);

Delay11No2_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_1_cast <= Delay11No2_out;
Delay5No14_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_2_cast <= Delay5No14_out;
   MUX_Add71_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No2_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay5No14_out_to_MUX_Add71_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add71_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add71_impl_0_out,
                 Y => Delay1No74_out);

SharedReg114_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg126_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_2_cast <= SharedReg126_out;
   MUX_Add71_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Add71_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add71_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add71_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add81_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add81_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add81_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add81_impl_out,
                 X => Delay1No76_out_to_Add81_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add81_impl_parent_implementedSystem_port_1_cast);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay1No76_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product112_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product112_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product112_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_impl_out,
                 X => Delay1No78_out_to_Product112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product112_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product112_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_0_out,
                 Y => Delay1No78_out);

SharedReg131_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product112_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product113_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product113_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product113_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_impl_out,
                 X => Delay1No80_out_to_Product113_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product113_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg63_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast <= SharedReg63_out;
   MUX_Product113_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product113_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_impl_0_out,
                 Y => Delay1No80_out);

SharedReg131_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg17_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
   MUX_Product113_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product113_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product101_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product101_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product101_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product101_impl_out,
                 X => Delay1No82_out_to_Product101_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product101_impl_parent_implementedSystem_port_1_cast);

Delay5No17_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast <= Delay5No17_out;
SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Product101_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No17_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product101_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product101_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product101_impl_0_out,
                 Y => Delay1No82_out);

SharedReg60_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Product101_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product101_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product101_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product101_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product121_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product121_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product121_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product121_impl_out,
                 X => Delay1No84_out_to_Product121_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product121_impl_parent_implementedSystem_port_1_cast);

SharedReg63_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg130_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product121_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product121_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product121_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product121_impl_0_out,
                 Y => Delay1No84_out);

SharedReg8_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg130_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product121_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product121_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product121_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product121_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product141_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product141_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product141_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product141_impl_out,
                 X => Delay1No86_out_to_Product141_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product141_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg130_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product141_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product141_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product141_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product141_impl_0_out,
                 Y => Delay1No86_out);

SharedReg13_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg130_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product141_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product141_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product141_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product141_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product151_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product151_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product151_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product151_impl_out,
                 X => Delay1No88_out_to_Product151_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product151_impl_parent_implementedSystem_port_1_cast);

SharedReg64_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_1_cast <= SharedReg64_out;
SharedReg67_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_2_cast <= SharedReg67_out;
   MUX_Product151_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg64_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg67_out_to_MUX_Product151_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product151_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product151_impl_0_out,
                 Y => Delay1No88_out);

SharedReg28_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Product151_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product151_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product151_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product151_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product171_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product171_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product171_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product171_impl_out,
                 X => Delay1No90_out_to_Product171_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product171_impl_parent_implementedSystem_port_1_cast);

Delay2No22_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast <= Delay2No22_out;
SharedReg130_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product171_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No22_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product171_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product171_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product171_impl_0_out,
                 Y => Delay1No90_out);

SharedReg18_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg130_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product171_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product171_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product171_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product171_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product181_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product181_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product181_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product181_impl_out,
                 X => Delay1No92_out_to_Product181_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product181_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product181_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product181_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product181_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_impl_0_out,
                 Y => Delay1No92_out);

SharedReg131_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product181_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product181_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product181_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product181_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product212_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product212_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product212_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product212_impl_out,
                 X => Delay1No94_out_to_Product212_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product212_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg69_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
   MUX_Product212_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product212_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product212_impl_0_out,
                 Y => Delay1No94_out);

SharedReg131_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg2_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast <= SharedReg2_out;
   MUX_Product212_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product212_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product212_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product221_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product221_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product221_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_impl_out,
                 X => Delay1No96_out_to_Product221_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product221_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg70_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast <= SharedReg70_out;
   MUX_Product221_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg70_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product221_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_0_out,
                 Y => Delay1No96_out);

SharedReg131_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg17_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
   MUX_Product221_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product221_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product241_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product241_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product241_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product241_impl_out,
                 X => Delay1No98_out_to_Product241_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product241_impl_parent_implementedSystem_port_1_cast);

SharedReg70_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg130_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product241_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product241_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_0_out,
                 Y => Delay1No98_out);

SharedReg23_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg130_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product241_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product241_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product251_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product251_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product251_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product251_impl_out,
                 X => Delay1No100_out_to_Product251_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product251_impl_parent_implementedSystem_port_1_cast);

Delay5No18_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_1_cast <= Delay5No18_out;
SharedReg130_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product251_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No18_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product251_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product251_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product251_impl_0_out,
                 Y => Delay1No100_out);

SharedReg59_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg130_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product251_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product251_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product251_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product251_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product261_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product261_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product261_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product261_impl_out,
                 X => Delay1No102_out_to_Product261_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product261_impl_parent_implementedSystem_port_1_cast);

Delay5No19_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_1_cast <= Delay5No19_out;
SharedReg130_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product261_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No19_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product261_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product261_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product261_impl_0_out,
                 Y => Delay1No102_out);

SharedReg61_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg130_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product261_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product261_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product261_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product261_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product271_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product271_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product271_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product271_impl_out,
                 X => Delay1No104_out_to_Product271_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product271_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product271_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product271_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product271_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product271_impl_0_out,
                 Y => Delay1No104_out);

SharedReg131_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product271_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product271_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product271_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product271_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product312_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product312_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product312_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_impl_out,
                 X => Delay1No106_out_to_Product312_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product312_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg76_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast <= SharedReg76_out;
   MUX_Product312_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product312_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_0_out,
                 Y => Delay1No106_out);

SharedReg131_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg22_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
   MUX_Product312_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product312_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product321_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product321_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product321_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_impl_out,
                 X => Delay1No108_out_to_Product321_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product321_impl_parent_implementedSystem_port_1_cast);

Delay6No13_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast <= Delay6No13_out;
SharedReg130_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product321_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No13_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product321_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_0_out,
                 Y => Delay1No108_out);

SharedReg59_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg130_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product321_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product321_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product361_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product361_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product361_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product361_impl_out,
                 X => Delay1No110_out_to_Product361_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product361_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg78_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
   MUX_Product361_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Product361_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product361_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product361_impl_0_out,
                 Y => Delay1No110_out);

SharedReg18_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg7_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_2_cast <= SharedReg7_out;
   MUX_Product361_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product361_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product361_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product361_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product401_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product401_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product401_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product401_impl_out,
                 X => Delay1No112_out_to_Product401_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product401_impl_parent_implementedSystem_port_1_cast);

SharedReg77_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_1_cast <= SharedReg77_out;
SharedReg130_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product401_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg77_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product401_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product401_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product401_impl_0_out,
                 Y => Delay1No112_out);

SharedReg8_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg130_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product401_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product401_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product401_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product401_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product412_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product412_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product412_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product412_impl_out,
                 X => Delay1No114_out_to_Product412_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product412_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product412_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product412_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product412_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product412_impl_0_out,
                 Y => Delay1No114_out);

SharedReg131_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product412_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product412_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product412_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product412_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product431_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product431_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product431_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product431_impl_out,
                 X => Delay1No116_out_to_Product431_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product431_impl_parent_implementedSystem_port_1_cast);

Delay5No20_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_1_cast <= Delay5No20_out;
SharedReg130_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product431_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No20_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product431_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product431_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_impl_0_out,
                 Y => Delay1No116_out);

SharedReg60_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg130_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product431_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product431_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product431_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product431_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product471_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product471_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product471_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product471_impl_out,
                 X => Delay1No118_out_to_Product471_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product471_impl_parent_implementedSystem_port_1_cast);

SharedReg97_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg82_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
   MUX_Product471_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product471_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product471_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product471_impl_0_out,
                 Y => Delay1No118_out);

SharedReg136_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg12_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_2_cast <= SharedReg12_out;
   MUX_Product471_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product471_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product471_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product471_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product481_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product481_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product481_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product481_impl_out,
                 X => Delay1No120_out_to_Product481_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product481_impl_parent_implementedSystem_port_1_cast);

SharedReg98_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg130_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product481_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product481_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product481_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_impl_0_out,
                 Y => Delay1No120_out);

SharedReg136_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg130_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product481_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product481_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product481_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product491_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product491_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product491_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product491_impl_out,
                 X => Delay1No122_out_to_Product491_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product491_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg130_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product491_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product491_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product491_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_impl_0_out,
                 Y => Delay1No122_out);

SharedReg60_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg130_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product491_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product491_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product491_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product491_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product512_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product512_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product512_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product512_impl_out,
                 X => Delay1No124_out_to_Product512_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product512_impl_parent_implementedSystem_port_1_cast);

SharedReg85_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg130_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product512_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product512_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product512_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_impl_0_out,
                 Y => Delay1No124_out);

SharedReg23_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg130_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product512_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product512_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product512_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product512_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product54_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product54_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product54_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product54_impl_out,
                 X => Delay1No126_out_to_Product54_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product54_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg81_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
   MUX_Product54_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product54_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_impl_0_out,
                 Y => Delay1No126_out);

SharedReg131_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg12_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast <= SharedReg12_out;
   MUX_Product54_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product54_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product55_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product55_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product55_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_impl_out,
                 X => Delay1No128_out_to_Product55_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product55_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg86_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast <= SharedReg86_out;
   MUX_Product55_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg86_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product55_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_0_out,
                 Y => Delay1No128_out);

SharedReg131_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg27_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Product55_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product55_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product57_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product57_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product57_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product57_impl_out,
                 X => Delay1No130_out_to_Product57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product57_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product57_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product57_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_impl_0_out,
                 Y => Delay1No130_out);

SharedReg131_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg130_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product57_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product57_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product59_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product59_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product59_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product59_impl_out,
                 X => Delay1No132_out_to_Product59_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product59_impl_parent_implementedSystem_port_1_cast);

Delay5No22_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast <= Delay5No22_out;
SharedReg130_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product59_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No22_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product59_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product59_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_impl_0_out,
                 Y => Delay1No132_out);

SharedReg59_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg130_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product59_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product59_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product59_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product61_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product61_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product61_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product61_impl_out,
                 X => Delay1No134_out_to_Product61_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product61_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg89_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_2_cast <= SharedReg89_out;
   MUX_Product61_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Product61_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product61_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_impl_0_out,
                 Y => Delay1No134_out);

SharedReg3_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg27_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Product61_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product61_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product61_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product63_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product63_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product63_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product63_impl_out,
                 X => Delay1No136_out_to_Product63_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product63_impl_parent_implementedSystem_port_1_cast);

SharedReg90_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg130_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product63_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product63_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product63_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_impl_0_out,
                 Y => Delay1No136_out);

SharedReg23_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg130_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product63_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product63_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product63_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product65_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product65_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product65_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product65_impl_out,
                 X => Delay1No138_out_to_Product65_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product65_impl_parent_implementedSystem_port_1_cast);

SharedReg93_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast <= SharedReg93_out;
SharedReg130_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product65_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg93_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product65_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product65_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product65_impl_0_out,
                 Y => Delay1No138_out);

SharedReg13_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg130_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product65_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product65_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product65_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product65_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product66_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product66_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product66_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product66_impl_out,
                 X => Delay1No140_out_to_Product66_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product66_impl_parent_implementedSystem_port_1_cast);

Delay5No23_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast <= Delay5No23_out;
SharedReg130_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product66_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No23_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product66_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product66_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_impl_0_out,
                 Y => Delay1No140_out);

SharedReg61_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg130_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product66_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product66_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product66_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product67_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product67_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product67_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product67_impl_out,
                 X => Delay1No142_out_to_Product67_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product67_impl_parent_implementedSystem_port_1_cast);

Delay6No15_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast <= Delay6No15_out;
SharedReg130_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product67_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No15_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product67_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_impl_0_out,
                 Y => Delay1No142_out);

SharedReg59_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg130_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product67_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product67_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Product68_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Product68_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Product68_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_impl_out,
                 X => Delay1No144_out_to_Product68_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Product68_impl_parent_implementedSystem_port_1_cast);

Delay6No16_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast <= Delay6No16_out;
SharedReg92_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast <= SharedReg92_out;
   MUX_Product68_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No16_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg92_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product68_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_impl_0_out,
                 Y => Delay1No144_out);

SharedReg60_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg2_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast <= SharedReg2_out;
   MUX_Product68_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product68_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product72_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product72_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product72_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product72_impl_out,
                 X => Delay1No146_out_to_Product72_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product72_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg15_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product72_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product72_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_0_out,
                 Y => Delay1No146_out);

SharedReg61_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg25_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Product72_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product72_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product73_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product73_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product73_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product73_impl_out,
                 X => Delay1No148_out_to_Product73_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product73_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg10_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Product73_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product73_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product73_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product73_impl_0_out,
                 Y => Delay1No148_out);

SharedReg24_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg25_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Product73_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product73_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product73_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product73_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product76_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product76_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product76_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product76_impl_out,
                 X => Delay1No150_out_to_Product76_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product76_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg130_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product76_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product76_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product76_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_impl_0_out,
                 Y => Delay1No150_out);

SharedReg61_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg130_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product76_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product76_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product76_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product77_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product77_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product77_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product77_impl_out,
                 X => Delay1No152_out_to_Product77_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product77_impl_parent_implementedSystem_port_1_cast);

SharedReg16_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg97_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast <= SharedReg97_out;
   MUX_Product77_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg97_out_to_MUX_Product77_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product77_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product77_impl_0_out,
                 Y => Delay1No152_out);

SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg132_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product77_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product77_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product77_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product77_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product81_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product81_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product81_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product81_impl_out,
                 X => Delay1No154_out_to_Product81_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product81_impl_parent_implementedSystem_port_1_cast);

Delay2No29_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast <= Delay2No29_out;
Delay11No_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast <= Delay11No_out;
   MUX_Product81_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No29_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No_out_to_MUX_Product81_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product81_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product81_impl_0_out,
                 Y => Delay1No154_out);

SharedReg133_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg62_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast <= SharedReg62_out;
   MUX_Product81_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Product81_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product81_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product81_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product82_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product82_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product82_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product82_impl_out,
                 X => Delay1No156_out_to_Product82_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product82_impl_parent_implementedSystem_port_1_cast);

SharedReg99_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg5_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Product82_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product82_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product82_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product82_impl_0_out,
                 Y => Delay1No156_out);

SharedReg136_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg20_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
   MUX_Product82_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product82_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product82_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product82_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product83_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product83_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product83_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product83_impl_out,
                 X => Delay1No158_out_to_Product83_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product83_impl_parent_implementedSystem_port_1_cast);

SharedReg100_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
   MUX_Product83_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Product83_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product83_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product83_impl_0_out,
                 Y => Delay1No158_out);

SharedReg133_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg20_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
   MUX_Product83_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product83_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product83_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product83_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product84_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product84_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product84_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product84_impl_out,
                 X => Delay1No160_out_to_Product84_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product84_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg5_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Product84_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product84_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product84_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product84_impl_0_out,
                 Y => Delay1No160_out);

SharedReg29_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
SharedReg25_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Product84_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product84_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product84_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product84_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product87_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product87_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product87_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product87_impl_out,
                 X => Delay1No162_out_to_Product87_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product87_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg99_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast <= SharedReg99_out;
   MUX_Product87_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg99_out_to_MUX_Product87_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product87_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product87_impl_0_out,
                 Y => Delay1No162_out);

SharedReg61_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg2_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast <= SharedReg2_out;
   MUX_Product87_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Product87_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product87_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product87_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product90_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product90_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product90_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product90_impl_out,
                 X => Delay1No164_out_to_Product90_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product90_impl_parent_implementedSystem_port_1_cast);

SharedReg104_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg102_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_2_cast <= SharedReg102_out;
   MUX_Product90_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Product90_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product90_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product90_impl_0_out,
                 Y => Delay1No164_out);

SharedReg136_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg132_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product90_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product90_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product90_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product90_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product91_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product91_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product91_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product91_impl_out,
                 X => Delay1No166_out_to_Product91_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product91_impl_parent_implementedSystem_port_1_cast);

SharedReg101_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg103_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_2_cast <= SharedReg103_out;
   MUX_Product91_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg103_out_to_MUX_Product91_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product91_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product91_impl_0_out,
                 Y => Delay1No166_out);

SharedReg137_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg132_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product91_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product91_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product91_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product91_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product93_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product93_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product93_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product93_impl_out,
                 X => Delay1No168_out_to_Product93_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product93_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg104_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_2_cast <= SharedReg104_out;
   MUX_Product93_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Product93_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product93_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product93_impl_0_out,
                 Y => Delay1No168_out);

SharedReg136_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg132_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product93_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product93_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product93_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product93_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product96_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product96_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product96_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product96_impl_out,
                 X => Delay1No170_out_to_Product96_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product96_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
   MUX_Product96_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Product96_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product96_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product96_impl_0_out,
                 Y => Delay1No170_out);

SharedReg19_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg10_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Product96_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product96_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product96_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product96_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product98_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product98_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product98_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product98_impl_out,
                 X => Delay1No172_out_to_Product98_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product98_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg25_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Product98_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product98_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product98_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product98_impl_0_out,
                 Y => Delay1No172_out);

SharedReg60_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg15_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product98_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product98_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product98_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product98_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product99_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product99_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product99_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product99_impl_out,
                 X => Delay1No174_out_to_Product99_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product99_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg110_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
   MUX_Product99_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Product99_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product99_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product99_impl_0_out,
                 Y => Delay1No174_out);

SharedReg60_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg132_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product99_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product99_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product99_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product99_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Subtract12_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_impl_out,
                 X => Delay1No176_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast);

SharedReg106_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
Delay10No11_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast <= Delay10No11_out;
   MUX_Subtract12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay10No11_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract12_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_0_out,
                 Y => Delay1No176_out);

Delay2No14_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast <= Delay2No14_out;
SharedReg42_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
   MUX_Subtract12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No14_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract12_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Subtract1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract1_impl_out,
                 X => Delay1No178_out_to_Subtract1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Subtract1_impl_parent_implementedSystem_port_1_cast);

Delay7No_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast <= Delay7No_out;
Delay2No18_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast <= Delay2No18_out;
   MUX_Subtract1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay2No18_out_to_MUX_Subtract1_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract1_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_impl_0_out,
                 Y => Delay1No178_out);

Delay2No15_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast <= Delay2No15_out;
SharedReg51_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg51_out;
   MUX_Subtract1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No15_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Subtract1_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract1_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Subtract2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_impl_out,
                 X => Delay1No180_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast);

SharedReg65_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
Delay2No23_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast <= Delay2No23_out;
   MUX_Subtract2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay2No23_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract2_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_0_out,
                 Y => Delay1No180_out);

SharedReg49_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg60_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg60_out;
   MUX_Subtract2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract2_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Subtract4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_impl_out,
                 X => Delay1No182_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast);

Delay11No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast <= Delay11No3_out;
Delay7No4_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast <= Delay7No4_out;
   MUX_Subtract4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No3_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay7No4_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract4_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_0_out,
                 Y => Delay1No182_out);

Delay2No16_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast <= Delay2No16_out;
SharedReg46_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg46_out;
   MUX_Subtract4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No16_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg46_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract4_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Subtract5_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Subtract5_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Subtract5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_impl_out,
                 X => Delay1No184_out_to_Subtract5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Subtract5_impl_parent_implementedSystem_port_1_cast);

SharedReg79_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg79_out;
Delay10No12_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_2_cast <= Delay10No12_out;
   MUX_Subtract5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay10No12_out_to_MUX_Subtract5_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract5_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_impl_0_out,
                 Y => Delay1No184_out);

Delay2No10_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_1_cast <= Delay2No10_out;
SharedReg48_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg48_out;
   MUX_Subtract5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No10_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Subtract5_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract5_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Subtract6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_impl_out,
                 X => Delay1No186_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay5No21_out,
                 Y => Delay1No186_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Subtract9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_impl_out,
                 X => Delay1No188_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay22No_out,
                 Y => Delay1No188_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Add32_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Add32_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Add32_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add32_impl_out,
                 X => Delay1No190_out_to_Add32_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Add32_impl_parent_implementedSystem_port_1_cast);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No461_out,
                 Y => Delay1No190_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay10No13_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Add11_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Add11_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Add11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_impl_out,
                 X => Delay1No192_out_to_Add11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Add11_impl_parent_implementedSystem_port_1_cast);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay61No_out,
                 Y => Delay1No192_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Add13_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Add13_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Add13_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add13_impl_out,
                 X => Delay1No194_out_to_Add13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Add13_impl_parent_implementedSystem_port_1_cast);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay79No_out,
                 Y => Delay1No194_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Add15_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Add15_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Add15_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_impl_out,
                 X => Delay1No196_out_to_Add15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Add15_impl_parent_implementedSystem_port_1_cast);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay81No_out,
                 Y => Delay1No196_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Add211_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Add211_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Add211_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add211_impl_out,
                 X => Delay1No198_out_to_Add211_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Add211_impl_parent_implementedSystem_port_1_cast);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay19No1_out,
                 Y => Delay1No198_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Add4_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Add4_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Add4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add4_impl_out,
                 X => Delay1No200_out_to_Add4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Add4_impl_parent_implementedSystem_port_1_cast);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay29No_out,
                 Y => Delay1No200_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Add6_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Add6_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Add6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_impl_out,
                 X => Delay1No202_out_to_Add6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Add6_impl_parent_implementedSystem_port_1_cast);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay31No_out,
                 Y => Delay1No202_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Add9_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Add9_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Add9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_impl_out,
                 X => Delay1No204_out_to_Add9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Add9_impl_parent_implementedSystem_port_1_cast);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay51No_out,
                 Y => Delay1No204_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => Delay1No205_out);
   Constant1_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_impl_out);

Delay1No206_out_to_Divide_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Divide_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Divide_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_impl_out,
                 X => Delay1No206_out_to_Divide_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Divide_impl_parent_implementedSystem_port_1_cast);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay107No_out,
                 Y => Delay1No206_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No412_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product115_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product115_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product115_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product115_impl_out,
                 X => Delay1No208_out_to_Product115_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product115_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg129_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast <= SharedReg129_out;
   MUX_Product115_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg129_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product115_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product115_impl_0_out,
                 Y => Delay1No208_out);

SharedReg19_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg134_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
   MUX_Product115_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product115_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product115_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product116_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product116_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product116_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product116_impl_out,
                 X => Delay1No210_out_to_Product116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product116_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg5_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Product116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product116_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_0_out,
                 Y => Delay1No210_out);

SharedReg136_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg25_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Product116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product116_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product10_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product10_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product10_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_impl_out,
                 X => Delay1No212_out_to_Product10_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product10_impl_parent_implementedSystem_port_1_cast);

Delay1No465_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast <= Delay1No465_out;
SharedReg20_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
   MUX_Product10_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay1No465_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product10_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_0_out,
                 Y => Delay1No212_out);

SharedReg136_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg15_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product10_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product10_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product11_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product11_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product11_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_impl_out,
                 X => Delay1No214_out_to_Product11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product11_impl_parent_implementedSystem_port_1_cast);

SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast <= SharedReg120_out;
SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg120_out;
   MUX_Product11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product11_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_0_out,
                 Y => Delay1No214_out);

SharedReg138_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg138_out;
SharedReg132_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg138_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product11_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product12_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product12_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product12_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_impl_out,
                 X => Delay1No216_out_to_Product12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product12_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg121_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_2_cast <= SharedReg121_out;
   MUX_Product12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Product12_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product12_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_impl_0_out,
                 Y => Delay1No216_out);

SharedReg60_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg134_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
   MUX_Product12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Product12_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product12_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product13_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product13_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product13_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_impl_out,
                 X => Delay1No218_out_to_Product13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product13_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
   MUX_Product13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product13_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_0_out,
                 Y => Delay1No218_out);

SharedReg136_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg10_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Product13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product13_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product14_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product14_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product14_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product14_impl_out,
                 X => Delay1No220_out_to_Product14_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product14_impl_parent_implementedSystem_port_1_cast);

SharedReg123_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast <= SharedReg123_out;
Delay1No322_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast <= Delay1No322_out;
   MUX_Product14_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No322_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product14_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_impl_0_out,
                 Y => Delay1No220_out);

SharedReg138_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast <= SharedReg138_out;
SharedReg130_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product14_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg138_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product14_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product15_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product15_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product15_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product15_impl_out,
                 X => Delay1No222_out_to_Product15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product15_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
Delay1No323_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast <= Delay1No323_out;
   MUX_Product15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No323_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product15_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product15_impl_0_out,
                 Y => Delay1No222_out);

SharedReg21_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg130_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product15_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product15_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product16_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product16_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product16_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product16_impl_out,
                 X => Delay1No224_out_to_Product16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product16_impl_parent_implementedSystem_port_1_cast);

SharedReg125_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg125_out;
Delay1No324_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast <= Delay1No324_out;
   MUX_Product16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No324_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product16_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_0_out,
                 Y => Delay1No224_out);

SharedReg133_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg130_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Product16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product16_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Product17_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Product17_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Product17_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_impl_out,
                 X => Delay1No226_out_to_Product17_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Product17_impl_parent_implementedSystem_port_1_cast);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => Delay1No226_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Product18_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Product18_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Product18_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_impl_out,
                 X => Delay1No228_out_to_Product18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Product18_impl_parent_implementedSystem_port_1_cast);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay1No228_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product19_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product19_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product19_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_impl_out,
                 X => Delay1No230_out_to_Product19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product19_impl_parent_implementedSystem_port_1_cast);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No440_out,
                 Y => Delay1No230_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product213_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product213_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product213_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_impl_out,
                 X => Delay1No232_out_to_Product213_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product213_impl_parent_implementedSystem_port_1_cast);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => Delay1No232_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product20_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product20_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product20_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product20_impl_out,
                 X => Delay1No234_out_to_Product20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product20_impl_parent_implementedSystem_port_1_cast);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No441_out,
                 Y => Delay1No234_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product21_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product21_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product21_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_impl_out,
                 X => Delay1No236_out_to_Product21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product21_impl_parent_implementedSystem_port_1_cast);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => Delay1No236_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Product22_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Product22_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Product22_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_impl_out,
                 X => Delay1No238_out_to_Product22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Product22_impl_parent_implementedSystem_port_1_cast);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No442_out,
                 Y => Delay1No238_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Product23_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Product23_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Product23_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_impl_out,
                 X => Delay1No240_out_to_Product23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Product23_impl_parent_implementedSystem_port_1_cast);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No443_out,
                 Y => Delay1No240_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product26_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product26_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product26_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_impl_out,
                 X => Delay1No242_out_to_Product26_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product26_impl_parent_implementedSystem_port_1_cast);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay2No39_out,
                 Y => Delay1No242_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product27_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product27_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product27_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_impl_out,
                 X => Delay1No244_out_to_Product27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product27_impl_parent_implementedSystem_port_1_cast);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay1No244_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product28_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product28_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product28_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_impl_out,
                 X => Delay1No246_out_to_Product28_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product28_impl_parent_implementedSystem_port_1_cast);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No445_out,
                 Y => Delay1No246_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product29_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product29_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product29_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product29_impl_out,
                 X => Delay1No248_out_to_Product29_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product29_impl_parent_implementedSystem_port_1_cast);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No446_out,
                 Y => Delay1No248_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Product3_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Product3_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Product3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product3_impl_out,
                 X => Delay1No250_out_to_Product3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Product3_impl_parent_implementedSystem_port_1_cast);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay1No250_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Product30_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Product30_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Product30_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product30_impl_out,
                 X => Delay1No252_out_to_Product30_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Product30_impl_parent_implementedSystem_port_1_cast);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay1No252_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product31_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product31_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product31_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_impl_out,
                 X => Delay1No254_out_to_Product31_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product31_impl_parent_implementedSystem_port_1_cast);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No448_out,
                 Y => Delay1No254_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product32_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product32_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product32_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_impl_out,
                 X => Delay1No256_out_to_Product32_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product32_impl_parent_implementedSystem_port_1_cast);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No449_out,
                 Y => Delay1No256_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product33_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product33_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product33_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_impl_out,
                 X => Delay1No258_out_to_Product33_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product33_impl_parent_implementedSystem_port_1_cast);

Delay1No450_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast <= Delay1No450_out;
SharedReg_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
   MUX_Product33_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay1No450_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product33_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_0_out,
                 Y => Delay1No258_out);

SharedReg135_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg15_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Product33_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product33_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product34_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product34_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product34_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product34_impl_out,
                 X => Delay1No260_out_to_Product34_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product34_impl_parent_implementedSystem_port_1_cast);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => Delay1No260_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Product36_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Product36_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Product36_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product36_impl_out,
                 X => Delay1No262_out_to_Product36_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Product36_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg5_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Product36_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product36_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_impl_0_out,
                 Y => Delay1No262_out);

SharedReg21_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg10_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Product36_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product36_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Product37_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Product37_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Product37_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_impl_out,
                 X => Delay1No264_out_to_Product37_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Product37_impl_parent_implementedSystem_port_1_cast);

SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast <= SharedReg128_out;
SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast <= SharedReg128_out;
   MUX_Product37_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product37_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_0_out,
                 Y => Delay1No264_out);

SharedReg133_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg132_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Product37_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product37_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product38_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product38_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product38_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_impl_out,
                 X => Delay1No266_out_to_Product38_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product38_impl_parent_implementedSystem_port_1_cast);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay1No266_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product4_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product4_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_impl_out,
                 X => Delay1No268_out_to_Product4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product4_impl_parent_implementedSystem_port_1_cast);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No447_out,
                 Y => Delay1No268_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Product43_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Product43_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Product43_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product43_impl_out,
                 X => Delay1No270_out_to_Product43_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Product43_impl_parent_implementedSystem_port_1_cast);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay2No41_out,
                 Y => Delay1No270_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Product44_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Product44_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Product44_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product44_impl_out,
                 X => Delay1No272_out_to_Product44_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Product44_impl_parent_implementedSystem_port_1_cast);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No456_out,
                 Y => Delay1No272_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Product45_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Product45_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Product45_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product45_impl_out,
                 X => Delay1No274_out_to_Product45_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Product45_impl_parent_implementedSystem_port_1_cast);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => Delay1No274_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Product46_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Product46_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Product46_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product46_impl_out,
                 X => Delay1No276_out_to_Product46_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Product46_impl_parent_implementedSystem_port_1_cast);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No457_out,
                 Y => Delay1No276_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product47_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product47_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product47_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product47_impl_out,
                 X => Delay1No278_out_to_Product47_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product47_impl_parent_implementedSystem_port_1_cast);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No458_out,
                 Y => Delay1No278_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product48_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product48_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product48_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product48_impl_out,
                 X => Delay1No280_out_to_Product48_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product48_impl_parent_implementedSystem_port_1_cast);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay1No280_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Product49_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Product49_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Product49_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product49_impl_out,
                 X => Delay1No282_out_to_Product49_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Product49_impl_parent_implementedSystem_port_1_cast);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No459_out,
                 Y => Delay1No282_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Product5_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Product5_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Product5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_impl_out,
                 X => Delay1No284_out_to_Product5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Product5_impl_parent_implementedSystem_port_1_cast);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No454_out,
                 Y => Delay1No284_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Product50_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Product50_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Product50_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_impl_out,
                 X => Delay1No286_out_to_Product50_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Product50_impl_parent_implementedSystem_port_1_cast);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No460_out,
                 Y => Delay1No286_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Product7_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Product7_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Product7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product7_impl_out,
                 X => Delay1No288_out_to_Product7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Product7_impl_parent_implementedSystem_port_1_cast);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay2No42_out,
                 Y => Delay1No288_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product8_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product8_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product8_impl_out,
                 X => Delay1No290_out_to_Product8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product8_impl_parent_implementedSystem_port_1_cast);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay1No464_out,
                 Y => Delay1No290_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product9_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product9_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product9_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_impl_out,
                 X => Delay1No292_out_to_Product9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product9_impl_parent_implementedSystem_port_1_cast);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => Delay1No292_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Subtract_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Subtract_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Subtract_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract_impl_out,
                 X => Delay1No294_out_to_Subtract_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Subtract_impl_parent_implementedSystem_port_1_cast);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Delay49No_out,
                 Y => Delay1No294_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => Delay1No295_out);
   Constant_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_impl_out);

   Delay5No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_out,
                 Y => Delay5No_out);

   Delay11No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => Delay11No_out);

   Delay5No7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_out,
                 Y => Delay5No7_out);

   Delay5No14_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_out,
                 Y => Delay5No14_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_out,
                 Y => Delay1No322_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_out,
                 Y => Delay1No323_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_out,
                 Y => Delay1No324_out);

   Delay92No_instance: Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=91 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => Delay92No_out);

   Delay2No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay2No10_out);

   Delay95No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => Delay95No_out);

   Delay97No_instance: Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=92 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => Delay97No_out);

   Delay97No1_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => Delay97No1_out);

   Delay2No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => Delay2No11_out);

   Delay2No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => Delay2No13_out);

   Delay75No_instance: Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=74 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => Delay75No_out);

   Delay2No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay2No14_out);

   Delay82No_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay82No_out);

   Delay2No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => Delay2No15_out);

   Delay83No_instance: Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=82 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => Delay83No_out);

   Delay97No2_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => Delay97No2_out);

   Delay97No3_instance: Delay_34_DelayLength_96_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=96 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay97No3_out);

   Delay97No4_instance: Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=95 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => Delay97No4_out);

   Delay2No16_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add81_impl_out,
                 Y => Delay2No16_out);

   Delay92No2_instance: Delay_34_DelayLength_90_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=90 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay92No2_out);

   Delay17No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => Delay17No_out);

   Delay5No16_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => Delay5No16_out);

   Delay2No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay2No17_out);

   Delay17No1_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => Delay17No1_out);

   Delay20No_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => Delay20No_out);

   Delay7No_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => Delay7No_out);

   Delay4No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => Delay4No_out);

   Delay4No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay4No1_out);

   Delay2No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => Delay2No18_out);

   Delay5No17_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => Delay5No17_out);

   Delay11No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => Delay11No1_out);

   Delay6No12_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay6No12_out);

   Delay2No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay2No22_out);

   Delay11No2_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => Delay11No2_out);

   Delay2No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => Delay2No23_out);

   Delay10No11_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => Delay10No11_out);

   Delay2No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => Delay2No24_out);

   Delay5No18_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => Delay5No18_out);

   Delay5No19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => Delay5No19_out);

   Delay17No2_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => Delay17No2_out);

   Delay11No3_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => Delay11No3_out);

   Delay5No20_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => Delay5No20_out);

   Delay6No13_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => Delay6No13_out);

   Delay9No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => Delay9No_out);

   Delay7No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => Delay7No2_out);

   Delay5No21_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => Delay5No21_out);

   Delay5No22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => Delay5No22_out);

   Delay5No23_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => Delay5No23_out);

   Delay7No3_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => Delay7No3_out);

   Delay7No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => Delay7No4_out);

   Delay6No15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay6No15_out);

   Delay6No16_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => Delay6No16_out);

   Delay17No3_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => Delay17No3_out);

   Delay10No12_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => Delay10No12_out);

   Delay2No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => Delay2No29_out);

   Delay25No_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => Delay25No_out);

   Delay19No_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => Delay19No_out);

   Delay22No_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => Delay22No_out);

   Delay15No_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => Delay15No_out);

   Delay9No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => Delay9No1_out);

   Delay12No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => Delay12No_out);

   Delay18No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => Delay18No_out);

   Delay11No4_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => Delay11No4_out);

   Delay2No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => Delay2No31_out);

   Delay2No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => Delay2No34_out);

   Delay2No36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_impl_out,
                 Y => Delay2No36_out);

   Delay2No38_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_impl_out,
                 Y => Delay2No38_out);

   Delay1No405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add32_impl_out,
                 Y => Delay1No405_out);

   Delay1No408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_impl_out,
                 Y => Delay1No408_out);

   Delay1No410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add13_impl_out,
                 Y => Delay1No410_out);

   Delay1No412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_impl_out,
                 Y => Delay1No412_out);

   Delay1No413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add211_impl_out,
                 Y => Delay1No413_out);

   Delay1No415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add4_impl_out,
                 Y => Delay1No415_out);

   Delay1No417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_impl_out,
                 Y => Delay1No417_out);

   Delay1No420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_impl_out,
                 Y => Delay1No420_out);

   Delay107No_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_impl_out,
                 Y => Delay107No_out);

   Delay66No_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => Delay66No_out);

   Delay61No_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => Delay61No_out);

   Delay64No_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_impl_out,
                 Y => Delay64No_out);

   Delay1No440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_impl_out,
                 Y => Delay1No440_out);

   Delay1No441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_impl_out,
                 Y => Delay1No441_out);

   Delay81No_instance: Delay_34_DelayLength_81_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=81 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_impl_out,
                 Y => Delay81No_out);

   Delay51No_instance: Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=51 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product20_impl_out,
                 Y => Delay51No_out);

   Delay1No442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_impl_out,
                 Y => Delay1No442_out);

   Delay1No443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_impl_out,
                 Y => Delay1No443_out);

   Delay46No_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_impl_out,
                 Y => Delay46No_out);

   Delay2No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => Delay2No39_out);

   Delay49No_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_impl_out,
                 Y => Delay49No_out);

   Delay1No445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_impl_out,
                 Y => Delay1No445_out);

   Delay1No446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_impl_out,
                 Y => Delay1No446_out);

   Delay36No_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product29_impl_out,
                 Y => Delay36No_out);

   Delay1No447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product3_impl_out,
                 Y => Delay1No447_out);

   Delay1No448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product30_impl_out,
                 Y => Delay1No448_out);

   Delay1No449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_impl_out,
                 Y => Delay1No449_out);

   Delay31No_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_impl_out,
                 Y => Delay31No_out);

   Delay1No450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product34_impl_out,
                 Y => Delay1No450_out);

   Delay34No_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => Delay34No_out);

   Delay29No_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_impl_out,
                 Y => Delay29No_out);

   Delay1No454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_impl_out,
                 Y => Delay1No454_out);

   Delay25No1_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => Delay25No1_out);

   Delay2No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => Delay2No41_out);

   Delay1No456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product43_impl_out,
                 Y => Delay1No456_out);

   Delay19No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product44_impl_out,
                 Y => Delay19No1_out);

   Delay1No457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product45_impl_out,
                 Y => Delay1No457_out);

   Delay1No458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product46_impl_out,
                 Y => Delay1No458_out);

   Delay14No_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product47_impl_out,
                 Y => Delay14No_out);

   Delay1No459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product48_impl_out,
                 Y => Delay1No459_out);

   Delay1No460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product49_impl_out,
                 Y => Delay1No460_out);

   Delay76No_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_impl_out,
                 Y => Delay76No_out);

   Delay1No461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_impl_out,
                 Y => Delay1No461_out);

   Delay10No13_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => Delay10No13_out);

   Delay2No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => Delay2No42_out);

   Delay1No464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product7_impl_out,
                 Y => Delay1No464_out);

   Delay79No_instance: Delay_34_DelayLength_79_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=79 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product8_impl_out,
                 Y => Delay79No_out);

   Delay1No465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_impl_out,
                 Y => Delay1No465_out);

   Delay1No466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract_impl_out,
                 Y => Delay1No466_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_impl_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_impl_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_impl_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_impl_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_impl_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_impl_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_impl_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_impl_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=92 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_impl_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_impl_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add151_impl_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_impl_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add19_impl_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add210_impl_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add20_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add21_impl_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_impl_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_impl_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add27_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add29_impl_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add31_impl_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add51_impl_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add61_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add71_impl_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_impl_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product101_impl_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product121_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product141_impl_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product151_impl_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product171_impl_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product181_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product212_impl_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product241_impl_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product251_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product261_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product271_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_impl_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product361_impl_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product401_impl_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product412_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product431_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product471_impl_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product481_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product491_impl_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product512_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product54_impl_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product57_impl_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product59_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product61_impl_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product63_impl_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product65_impl_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product66_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product67_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product72_impl_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product73_impl_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product76_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product77_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product81_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product82_impl_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product83_impl_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product84_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product87_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product90_impl_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product91_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product93_impl_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product96_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product98_impl_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product99_impl_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_impl_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract1_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_impl_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_impl_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product115_impl_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product116_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_impl_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_impl_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product14_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product15_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product16_impl_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product36_impl_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_impl_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);
end architecture;

