--------------------------------------------------------------------------------
--                         ModuloCounter_59_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_59_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_59_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 58 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_31_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_31_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_31_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_28_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_28_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_28_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n352_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n352_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n352_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011101100000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n432_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n432_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n432_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011110110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n500_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n500_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n500_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011111110100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n532_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n532_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n532_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111100000001010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n129_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n129_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n129_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011000000010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_158_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_158_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_158_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111011000111100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_526_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_526_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_526_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100000000111000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_964_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_964_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_964_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100011100010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n529_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n529_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n529_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111100000001000100000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n464_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n464_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n464_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_29_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_29_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_29_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n336_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n336_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n336_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011101010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_3136_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_3136_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_3136_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101010001000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_3648_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_3648_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_3648_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101011001000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4110_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4110_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4110_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100000000111000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4478_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4478_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4478_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100010111111000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4737_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4737_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4737_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100101000000100000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4868_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4868_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4868_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100110000010000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_22_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_22_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_22_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001101100000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_1472_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1472_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1472_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100101110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_2008_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_2008_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_2008_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100111110110000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_2576_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_2576_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_2576_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101001000010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_8_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_8_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_8_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n17_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n17_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n17_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111001100010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n59_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n59_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n59_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111010011011000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n116_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n116_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n116_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111010111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n188_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n188_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n188_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011001111000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n268_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n268_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n268_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011100001100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid317669
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid317669 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid317669 is
signal XX_m317670 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m317670 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m317670 <= X ;
   YY_m317670 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid317673
--                   (IntAdderClassical_33_f500_uid317675)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid317673 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid317673 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid317669 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid317673 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid317669  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid317673  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_56_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_56_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_56_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_36_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_36_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_36_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_50_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_50_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_50_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_26_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_26_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_26_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
         iS_19 when "10011",
         iS_20 when "10100",
         iS_21 when "10101",
         iS_22 when "10110",
         iS_23 when "10111",
         iS_24 when "11000",
         iS_25 when "11001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_11_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_11_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_11_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid317796_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid317798)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid317796_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid317796_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid317801
--                  (IntAdderAlternative_27_f250_uid317805)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid317801 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid317801 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid317808
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid317808 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid317808 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid317811
--                   (IntAdderClassical_34_f250_uid317813)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid317811 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid317811 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid317796
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid317796 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid317796 is
   component FPAdd_8_23_uid317796_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid317801 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid317808 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid317811 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid317796_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid317801  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid317808  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid317811  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid317796 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid317796  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_59_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_59_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_59_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      Y <= s32;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 52 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      Y <= s51;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      Y <= s37;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 70 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      Y <= s69;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_160_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 160 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_160_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_160_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
signal s154 : std_logic_vector(33 downto 0) := (others => '0');
signal s155 : std_logic_vector(33 downto 0) := (others => '0');
signal s156 : std_logic_vector(33 downto 0) := (others => '0');
signal s157 : std_logic_vector(33 downto 0) := (others => '0');
signal s158 : std_logic_vector(33 downto 0) := (others => '0');
signal s159 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
      s154 <= "0000000000000000000000000000000000";
      s155 <= "0000000000000000000000000000000000";
      s156 <= "0000000000000000000000000000000000";
      s157 <= "0000000000000000000000000000000000";
      s158 <= "0000000000000000000000000000000000";
      s159 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      s154 <= s153;
      s155 <= s154;
      s156 <= s155;
      s157 <= s156;
      s158 <= s157;
      s159 <= s158;
      Y <= s159;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 105 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      Y <= s104;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 146 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      Y <= s145;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 103 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      Y <= s102;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 48 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      Y <= s47;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 66 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      Y <= s65;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_101_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 101 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_101_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_101_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      Y <= s100;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 115 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      Y <= s114;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_154_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 154 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_154_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_154_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
signal s147 : std_logic_vector(33 downto 0) := (others => '0');
signal s148 : std_logic_vector(33 downto 0) := (others => '0');
signal s149 : std_logic_vector(33 downto 0) := (others => '0');
signal s150 : std_logic_vector(33 downto 0) := (others => '0');
signal s151 : std_logic_vector(33 downto 0) := (others => '0');
signal s152 : std_logic_vector(33 downto 0) := (others => '0');
signal s153 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
      s147 <= "0000000000000000000000000000000000";
      s148 <= "0000000000000000000000000000000000";
      s149 <= "0000000000000000000000000000000000";
      s150 <= "0000000000000000000000000000000000";
      s151 <= "0000000000000000000000000000000000";
      s152 <= "0000000000000000000000000000000000";
      s153 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      s147 <= s146;
      s148 <= s147;
      s149 <= s148;
      s150 <= s149;
      s151 <= s150;
      s152 <= s151;
      s153 <= s152;
      Y <= s153;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "101010" when "000000",
      "100010" when "000001",
      "001010" when "000010",
      "001101" when "000011",
      "001011" when "000100",
      "010100" when "000101",
      "000100" when "000110",
      "010111" when "000111",
      "100110" when "001000",
      "000000" when "001001",
      "000010" when "001010",
      "100001" when "001011",
      "101001" when "001100",
      "000101" when "001101",
      "011010" when "001110",
      "000001" when "001111",
      "000000" when "010000",
      "011110" when "010001",
      "000011" when "010010",
      "101000" when "010011",
      "011000" when "010100",
      "101101" when "010101",
      "101110" when "010110",
      "011011" when "010111",
      "000110" when "011000",
      "010011" when "011001",
      "101111" when "011010",
      "010101" when "011011",
      "100100" when "011100",
      "110011" when "011101",
      "100011" when "011110",
      "000000" when "011111",
      "000111" when "100000",
      "010001" when "100001",
      "110000" when "100010",
      "010000" when "100011",
      "110001" when "100100",
      "110110" when "100101",
      "010110" when "100110",
      "110111" when "100111",
      "011101" when "101000",
      "001000" when "101001",
      "011001" when "101010",
      "001100" when "101011",
      "101100" when "101100",
      "110101" when "101101",
      "100111" when "101110",
      "011100" when "101111",
      "110010" when "110000",
      "000000" when "110001",
      "001001" when "110010",
      "001111" when "110011",
      "100101" when "110100",
      "110100" when "110101",
      "100000" when "110110",
      "001110" when "110111",
      "011111" when "111000",
      "101011" when "111001",
      "010010" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100011" when "000000",
      "100100" when "000001",
      "001000" when "000010",
      "010000" when "000011",
      "001001" when "000100",
      "100001" when "000101",
      "100111" when "000110",
      "001100" when "000111",
      "101010" when "001000",
      "110011" when "001001",
      "110101" when "001010",
      "100000" when "001011",
      "000001" when "001100",
      "101100" when "001101",
      "110110" when "001110",
      "110100" when "001111",
      "000000" when "010000",
      "011101" when "010001",
      "100110" when "010010",
      "000000" when "010011",
      "001101" when "010100",
      "000010" when "010101",
      "000011" when "010110",
      "110111" when "010111",
      "101101" when "011000",
      "011001" when "011001",
      "000100" when "011010",
      "100010" when "011011",
      "101000" when "011100",
      "000110" when "011101",
      "100101" when "011110",
      "000000" when "011111",
      "101110" when "100000",
      "010111" when "100001",
      "000101" when "100010",
      "010011" when "100011",
      "110001" when "100100",
      "010101" when "100101",
      "001011" when "100110",
      "010110" when "100111",
      "011100" when "101000",
      "101111" when "101001",
      "001110" when "101010",
      "001010" when "101011",
      "011011" when "101100",
      "010100" when "101101",
      "101011" when "101110",
      "001111" when "101111",
      "110010" when "110000",
      "000000" when "110001",
      "110000" when "110010",
      "010010" when "110011",
      "101001" when "110100",
      "000111" when "110101",
      "011111" when "110110",
      "010001" when "110111",
      "011110" when "111000",
      "011010" when "111001",
      "011000" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001101" when "000000",
      "010111" when "000001",
      "010011" when "000010",
      "000000" when "000011",
      "000110" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "000010" when "000111",
      "000000" when "001000",
      "000001" when "001001",
      "011001" when "001010",
      "000000" when "001011",
      "010000" when "001100",
      "000011" when "001101",
      "001111" when "001110",
      "010110" when "001111",
      "000000" when "010000",
      "011000" when "010001",
      "000000" when "010010",
      "011010" when "010011",
      "001011" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "000000" when "010111",
      "000111" when "011000",
      "000000" when "011001",
      "000000" when "011010",
      "011101" when "011011",
      "011011" when "011100",
      "011100" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "001000" when "100000",
      "001001" when "100001",
      "000000" when "100010",
      "000000" when "100011",
      "011111" when "100100",
      "001010" when "100101",
      "001100" when "100110",
      "100000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "000000" when "101010",
      "011110" when "101011",
      "000100" when "101100",
      "000000" when "101101",
      "100010" when "101110",
      "100011" when "101111",
      "010101" when "110000",
      "000000" when "110001",
      "010100" when "110010",
      "010001" when "110011",
      "000101" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "010010" when "110111",
      "100001" when "111000",
      "000000" when "111001",
      "001110" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001000" when "000000",
      "010111" when "000001",
      "010100" when "000010",
      "000000" when "000011",
      "011100" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "100001" when "000111",
      "000000" when "001000",
      "100000" when "001001",
      "010010" when "001010",
      "000000" when "001011",
      "100011" when "001100",
      "100010" when "001101",
      "001010" when "001110",
      "000001" when "001111",
      "000000" when "010000",
      "011000" when "010001",
      "011111" when "010010",
      "000010" when "010011",
      "010101" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "000000" when "010111",
      "000111" when "011000",
      "000000" when "011001",
      "000000" when "011010",
      "000101" when "011011",
      "000011" when "011100",
      "000100" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "001111" when "100000",
      "010000" when "100001",
      "000000" when "100010",
      "000000" when "100011",
      "011101" when "100100",
      "010001" when "100101",
      "010110" when "100110",
      "011110" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "000000" when "101010",
      "000110" when "101011",
      "011001" when "101100",
      "000000" when "101101",
      "001101" when "101110",
      "001110" when "101111",
      "011011" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "001011" when "110011",
      "011010" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "010011" when "110111",
      "001100" when "111000",
      "000000" when "111001",
      "001001" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100100" when "000000",
      "001011" when "000001",
      "011000" when "000010",
      "011111" when "000011",
      "001111" when "000100",
      "010001" when "000101",
      "000000" when "000110",
      "100001" when "000111",
      "001110" when "001000",
      "000010" when "001001",
      "010110" when "001010",
      "100110" when "001011",
      "010100" when "001100",
      "000001" when "001101",
      "010111" when "001110",
      "010101" when "001111",
      "000000" when "010000",
      "011101" when "010001",
      "101001" when "010010",
      "011010" when "010011",
      "101100" when "010100",
      "101011" when "010101",
      "000000" when "010110",
      "000100" when "010111",
      "000110" when "011000",
      "000000" when "011001",
      "100000" when "011010",
      "010010" when "011011",
      "011011" when "011100",
      "101101" when "011101",
      "101110" when "011110",
      "000000" when "011111",
      "000111" when "100000",
      "101111" when "100001",
      "110001" when "100010",
      "000000" when "100011",
      "100010" when "100100",
      "010011" when "100101",
      "001001" when "100110",
      "101000" when "100111",
      "011100" when "101000",
      "000000" when "101001",
      "100111" when "101010",
      "000000" when "101011",
      "101010" when "101100",
      "010000" when "101101",
      "100101" when "101110",
      "011001" when "101111",
      "110000" when "110000",
      "000000" when "110001",
      "011110" when "110010",
      "001010" when "110011",
      "100011" when "110100",
      "000000" when "110101",
      "001100" when "110110",
      "001000" when "110111",
      "000011" when "111000",
      "000101" when "111001",
      "001101" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011111" when "000000",
      "010001" when "000001",
      "001111" when "000010",
      "100111" when "000011",
      "010101" when "000100",
      "011100" when "000101",
      "000000" when "000110",
      "000000" when "000111",
      "010100" when "001000",
      "101110" when "001001",
      "110000" when "001010",
      "100001" when "001011",
      "001110" when "001100",
      "101101" when "001101",
      "110001" when "001110",
      "101111" when "001111",
      "000000" when "010000",
      "100010" when "010001",
      "000001" when "010010",
      "011001" when "010011",
      "000100" when "010100",
      "000011" when "010101",
      "000000" when "010110",
      "100101" when "010111",
      "101010" when "011000",
      "000000" when "011001",
      "101000" when "011010",
      "001100" when "011011",
      "011010" when "011100",
      "000101" when "011101",
      "000110" when "011110",
      "000000" when "011111",
      "101011" when "100000",
      "000111" when "100001",
      "001001" when "100010",
      "000000" when "100011",
      "011101" when "100100",
      "001101" when "100101",
      "001010" when "100110",
      "011000" when "100111",
      "011011" when "101000",
      "000000" when "101001",
      "010111" when "101010",
      "100011" when "101011",
      "000010" when "101100",
      "010110" when "101101",
      "100000" when "101110",
      "010000" when "101111",
      "001000" when "110000",
      "000000" when "110001",
      "100110" when "110010",
      "001011" when "110011",
      "011110" when "110100",
      "000000" when "110101",
      "010010" when "110110",
      "101100" when "110111",
      "100100" when "111000",
      "101001" when "111001",
      "010011" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00110" when "000000",
      "10101" when "000001",
      "00011" when "000010",
      "00000" when "000011",
      "01100" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "00010" when "000111",
      "00000" when "001000",
      "00001" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00000" when "001100",
      "01011" when "001101",
      "10000" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "10100" when "010001",
      "00000" when "010010",
      "10011" when "010011",
      "10001" when "010100",
      "00000" when "010101",
      "00000" when "010110",
      "00000" when "010111",
      "10111" when "011000",
      "00000" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00111" when "011100",
      "11001" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "00100" when "100000",
      "10010" when "100001",
      "00000" when "100010",
      "00000" when "100011",
      "00101" when "100100",
      "01000" when "100101",
      "00000" when "100110",
      "00000" when "100111",
      "00000" when "101000",
      "00000" when "101001",
      "00000" when "101010",
      "11000" when "101011",
      "01101" when "101100",
      "00000" when "101101",
      "01110" when "101110",
      "00000" when "101111",
      "00000" when "110000",
      "00000" when "110001",
      "00000" when "110010",
      "00000" when "110011",
      "10110" when "110100",
      "00000" when "110101",
      "00000" when "110110",
      "01010" when "110111",
      "01111" when "111000",
      "00000" when "111001",
      "01001" when "111010",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00110" when "000000",
      "10000" when "000001",
      "01001" when "000010",
      "00000" when "000011",
      "01101" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "11001" when "000111",
      "00000" when "001000",
      "11000" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00000" when "001100",
      "01100" when "001101",
      "10011" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "00010" when "010001",
      "10111" when "010010",
      "00001" when "010011",
      "10100" when "010100",
      "00000" when "010101",
      "00000" when "010110",
      "00000" when "010111",
      "00011" when "011000",
      "00000" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00111" when "011100",
      "00100" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "01111" when "100000",
      "10101" when "100001",
      "00000" when "100010",
      "00000" when "100011",
      "00101" when "100100",
      "01000" when "100101",
      "00000" when "100110",
      "00000" when "100111",
      "00000" when "101000",
      "00000" when "101001",
      "00000" when "101010",
      "10110" when "101011",
      "00000" when "101100",
      "00000" when "101101",
      "01110" when "101110",
      "00000" when "101111",
      "00000" when "110000",
      "00000" when "110001",
      "00000" when "110010",
      "00000" when "110011",
      "10001" when "110100",
      "00000" when "110101",
      "00000" when "110110",
      "01011" when "110111",
      "10010" when "111000",
      "00000" when "111001",
      "01010" when "111010",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0111" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0110" when "000111",
      "0000" when "001000",
      "0100" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "0001" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "1000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "1001" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "1010" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "0000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0010" when "110111",
      "0011" when "111000",
      "0000" when "111001",
      "0101" when "111010",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "0011" when "000000",
      "0000" when "000001",
      "0000" when "000010",
      "0000" when "000011",
      "0000" when "000100",
      "0000" when "000101",
      "0000" when "000110",
      "0101" when "000111",
      "0000" when "001000",
      "0110" when "001001",
      "0000" when "001010",
      "0000" when "001011",
      "0000" when "001100",
      "0000" when "001101",
      "0000" when "001110",
      "0000" when "001111",
      "0000" when "010000",
      "0000" when "010001",
      "0000" when "010010",
      "0000" when "010011",
      "1001" when "010100",
      "0000" when "010101",
      "0000" when "010110",
      "0000" when "010111",
      "0000" when "011000",
      "0000" when "011001",
      "0000" when "011010",
      "0000" when "011011",
      "0000" when "011100",
      "0000" when "011101",
      "0000" when "011110",
      "0000" when "011111",
      "0001" when "100000",
      "0000" when "100001",
      "0000" when "100010",
      "0000" when "100011",
      "0000" when "100100",
      "1010" when "100101",
      "0000" when "100110",
      "0000" when "100111",
      "0000" when "101000",
      "0000" when "101001",
      "0000" when "101010",
      "1000" when "101011",
      "0000" when "101100",
      "0000" when "101101",
      "0000" when "101110",
      "0000" when "101111",
      "0000" when "110000",
      "0000" when "110001",
      "0000" when "110010",
      "0000" when "110011",
      "0000" when "110100",
      "0000" when "110101",
      "0000" when "110110",
      "0010" when "110111",
      "0100" when "111000",
      "0000" when "111001",
      "0111" when "111010",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 60 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      Y <= s59;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 40 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      Y <= s39;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 88 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      Y <= s87;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      Y <= s40;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 54 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      Y <= s53;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      Y <= s55;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 74 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      Y <= s73;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 86 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      Y <= s85;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 117 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      Y <= s116;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 59 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      Y <= s58;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_141_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 141 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_141_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_141_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      Y <= s140;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 50 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      Y <= s49;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      Y <= s62;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 82 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      Y <= s81;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          X_0 : in std_logic_vector(31 downto 0);
          X_1 : in std_logic_vector(31 downto 0);
          X_2 : in std_logic_vector(31 downto 0);
          X_3 : in std_logic_vector(31 downto 0);
          X_4 : in std_logic_vector(31 downto 0);
          X_5 : in std_logic_vector(31 downto 0);
          Y_0 : out std_logic_vector(31 downto 0);
          Y_1 : out std_logic_vector(31 downto 0);
          Y_2 : out std_logic_vector(31 downto 0);
          Y_3 : out std_logic_vector(31 downto 0);
          Y_4 : out std_logic_vector(31 downto 0);
          Y_5 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_59_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_31_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_28_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n352_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n432_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n500_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n532_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n129_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_158_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_526_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_964_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n529_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n464_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_29_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n336_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_3136_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_3648_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4110_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4478_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4737_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4868_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_22_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1472_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_2008_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_2576_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_8_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n17_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n59_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n116_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n188_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n268_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_56_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_36_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_50_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_26_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_11_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_59_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_160_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_101_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_154_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_141_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount591_out : std_logic_vector(5 downto 0) := (others => '0');
signal X_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant19_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant20_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant24_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant25_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant29_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant34_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product1_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum11_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum11_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum11_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay546No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay590No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay591No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay597No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay603No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay607No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay101No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay138No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay109No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay169No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay322No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay323No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay161No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay211No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay278No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay38No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay52No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay249No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay296No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay339No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay358No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay351No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay122No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay225No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay135No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay266No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay288No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay134No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_0_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_2_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_2_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_3_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_3_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product1_2_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product1_2_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay101No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay107No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay138No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No3_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay65No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay322No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay323No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay278No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay52No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay266No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay288No_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay109No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay161No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay91No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay211No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No2_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay38No_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay75No3_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay225No_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay135No3_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay13No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay169No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay122No1_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay590No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay591No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay597No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay603No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay546No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay134No1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay249No1_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay358No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay339No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay607No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Sum11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Sum11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Sum11_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Sum11_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay296No_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay351No2_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Y_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount591_instance: ModuloCounter_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount591_out);
X_0_IEEE <= X_0;
   X_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_0_out,
                 X => X_0_IEEE);
X_1_IEEE <= X_1;
   X_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_1_out,
                 X => X_1_IEEE);
X_2_IEEE <= X_2;
   X_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_2_out,
                 X => X_2_IEEE);
X_3_IEEE <= X_3;
   X_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_3_out,
                 X => X_3_IEEE);
X_4_IEEE <= X_4;
   X_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_4_out,
                 X => X_4_IEEE);
X_5_IEEE <= X_5;
   X_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_5_out,
                 X => X_5_IEEE);
   Constant_0_impl_instance: Constant_float_8_23_31_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_28_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);
   Constant10_0_impl_instance: Constant_float_8_23_n352_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant10_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_n432_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant12_0_impl_instance: Constant_float_8_23_n500_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant12_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_n532_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_n129_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_158_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_526_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_964_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_n529_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant19_0_impl_instance: Constant_float_8_23_n464_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant19_0_impl_out);
   Constant2_0_impl_instance: Constant_float_8_23_29_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant20_0_impl_instance: Constant_float_8_23_n336_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant20_0_impl_out);
   Constant21_0_impl_instance: Constant_float_8_23_3136_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant21_0_impl_out);
   Constant22_0_impl_instance: Constant_float_8_23_3648_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant22_0_impl_out);
   Constant23_0_impl_instance: Constant_float_8_23_4110_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant23_0_impl_out);
   Constant24_0_impl_instance: Constant_float_8_23_4478_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant24_0_impl_out);
   Constant25_0_impl_instance: Constant_float_8_23_4737_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant25_0_impl_out);
   Constant29_0_impl_instance: Constant_float_8_23_4868_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant29_0_impl_out);
   Constant3_0_impl_instance: Constant_float_8_23_22_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant3_0_impl_out);
   Constant32_0_impl_instance: Constant_float_8_23_1472_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant32_0_impl_out);
   Constant33_0_impl_instance: Constant_float_8_23_2008_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant33_0_impl_out);
   Constant34_0_impl_instance: Constant_float_8_23_2576_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant34_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_8_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_n17_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_n59_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_n116_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_n188_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_n268_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);

Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_0_impl_out,
                 X => Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast);

SharedReg339_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg339_out;
SharedReg341_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg343_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
SharedReg348_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg348_out;
SharedReg347_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg347_out;
SharedReg352_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg352_out;
Delay77No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast <= Delay77No1_out;
SharedReg353_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg353_out;
SharedReg354_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg354_out;
SharedReg358_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg358_out;
SharedReg365_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg365_out;
SharedReg366_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg366_out;
Delay101No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast <= Delay101No_out;
SharedReg369_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg369_out;
SharedReg368_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg368_out;
Delay107No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast <= Delay107No_out;
SharedReg371_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg371_out;
Delay91No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast <= Delay91No2_out;
SharedReg379_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg379_out;
Delay138No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast <= Delay138No_out;
SharedReg384_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg384_out;
SharedReg382_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg382_out;
SharedReg387_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg387_out;
SharedReg390_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg390_out;
SharedReg396_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg396_out;
SharedReg393_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg393_out;
SharedReg400_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg400_out;
Delay19No3_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast <= Delay19No3_out;
SharedReg404_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg404_out;
SharedReg410_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg410_out;
SharedReg409_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg409_out;
SharedReg415_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg415_out;
SharedReg420_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg420_out;
Delay65No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast <= Delay65No1_out;
SharedReg424_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg424_out;
Delay322No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast <= Delay322No1_out;
Delay323No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast <= Delay323No2_out;
SharedReg426_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg426_out;
SharedReg431_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg431_out;
SharedReg434_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg434_out;
SharedReg440_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg440_out;
SharedReg437_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg437_out;
SharedReg444_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg444_out;
SharedReg455_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg455_out;
Delay278No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast <= Delay278No_out;
SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg457_out;
SharedReg461_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg461_out;
SharedReg464_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg464_out;
SharedReg467_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg467_out;
SharedReg470_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg470_out;
SharedReg471_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg471_out;
Delay52No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast <= Delay52No2_out;
SharedReg476_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg476_out;
SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg475_out;
SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg475_out;
   MUX_Product_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg339_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg365_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg366_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay101No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg369_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg368_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay107No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg371_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay91No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg379_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay138No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg343_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg384_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg382_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg387_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg390_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg396_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg393_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg400_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay19No3_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg404_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg410_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg348_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg409_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg415_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg420_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay65No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg424_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => Delay322No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => Delay323No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg426_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg431_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg434_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg347_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg440_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg437_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg444_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg455_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay278No_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg457_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg461_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg464_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg467_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg352_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg470_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg471_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => Delay52No2_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg476_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg475_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => Delay77No1_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg353_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg354_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg358_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_0_impl_0_LUT_out,
                 oMux => MUX_Product_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg659_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg659_out;
SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg633_out;
SharedReg729_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg614_out;
SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg608_out;
SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg608_out;
SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg673_out;
SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg617_out;
SharedReg697_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg697_out;
SharedReg693_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg693_out;
SharedReg615_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg615_out;
SharedReg644_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg644_out;
SharedReg626_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg626_out;
SharedReg712_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg712_out;
SharedReg722_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg722_out;
SharedReg619_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg619_out;
SharedReg613_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg613_out;
SharedReg650_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg650_out;
SharedReg690_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg690_out;
SharedReg699_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg699_out;
SharedReg708_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg708_out;
SharedReg654_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg654_out;
SharedReg718_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg718_out;
SharedReg624_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg624_out;
SharedReg652_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg652_out;
SharedReg629_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg629_out;
SharedReg726_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg726_out;
SharedReg630_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg630_out;
SharedReg641_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg641_out;
SharedReg700_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg700_out;
SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg609_out;
SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg713_out;
SharedReg627_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg627_out;
SharedReg679_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg679_out;
SharedReg623_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg623_out;
SharedReg631_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg631_out;
Delay266No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast <= Delay266No1_out;
SharedReg618_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg618_out;
SharedReg728_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg728_out;
Delay288No_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast <= Delay288No_out;
SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg633_out;
SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg609_out;
SharedReg648_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg648_out;
SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg614_out;
SharedReg723_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg723_out;
SharedReg711_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg711_out;
SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg673_out;
SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg617_out;
SharedReg703_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg703_out;
SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg713_out;
SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg608_out;
SharedReg611_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg611_out;
SharedReg634_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg634_out;
SharedReg704_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg704_out;
SharedReg653_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg653_out;
   MUX_Product_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg659_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg693_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg615_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg644_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg626_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg712_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg722_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg619_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg613_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg650_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg690_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg699_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg708_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg654_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg718_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg624_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg652_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg629_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg726_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg630_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg641_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg729_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg700_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg627_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg679_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg623_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg631_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => Delay266No1_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg618_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg728_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => Delay288No_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg633_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg609_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg648_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg614_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg723_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg711_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg703_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg713_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg611_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg634_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg704_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg653_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg608_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg673_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg617_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg697_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_0_impl_1_LUT_out,
                 oMux => MUX_Product_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_2_impl_out,
                 X => Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast);

Delay18No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast <= Delay18No_out;
SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg340_out;
SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg340_out;
SharedReg346_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg346_out;
Delay102No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast <= Delay102No_out;
SharedReg350_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg350_out;
SharedReg360_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg360_out;
SharedReg362_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg373_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg373_out;
SharedReg372_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg372_out;
SharedReg377_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg377_out;
SharedReg386_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg386_out;
SharedReg383_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg383_out;
SharedReg388_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg388_out;
Delay111No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast <= Delay111No_out;
SharedReg395_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg395_out;
SharedReg399_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg399_out;
Delay109No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast <= Delay109No_out;
SharedReg406_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg406_out;
SharedReg419_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg419_out;
SharedReg418_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg418_out;
Delay161No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast <= Delay161No_out;
SharedReg439_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg439_out;
SharedReg449_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg449_out;
SharedReg446_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg446_out;
SharedReg451_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg451_out;
Delay76No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast <= Delay76No1_out;
SharedReg463_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg463_out;
SharedReg462_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg462_out;
SharedReg459_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg459_out;
SharedReg466_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg466_out;
Delay95No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast <= Delay95No_out;
SharedReg468_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg468_out;
Delay55No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast <= Delay55No1_out;
SharedReg476_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg476_out;
SharedReg477_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg477_out;
   MUX_Product_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_36_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay18No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg377_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg386_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg383_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg388_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay111No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg395_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg399_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay109No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg406_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg419_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg340_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg418_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay161No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg439_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg449_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg446_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg451_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay76No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg463_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg462_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg459_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg346_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg466_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => Delay95No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg468_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay55No1_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg476_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg477_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_4 => Delay102No_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg360_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg373_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg372_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_2_impl_0_LUT_out,
                 oMux => MUX_Product_2_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_0_out,
                 Y => Delay1No2_out);

SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg633_out;
SharedReg674_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg674_out;
SharedReg720_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg720_out;
SharedReg636_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg658_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg658_out;
SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg654_out;
SharedReg716_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg716_out;
SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg657_out;
SharedReg691_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg691_out;
SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg651_out;
SharedReg685_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg685_out;
SharedReg671_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg671_out;
SharedReg719_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg719_out;
SharedReg665_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg665_out;
SharedReg737_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg737_out;
SharedReg614_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg614_out;
SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg657_out;
SharedReg681_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg681_out;
SharedReg677_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg677_out;
SharedReg646_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg646_out;
SharedReg611_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg611_out;
SharedReg666_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg666_out;
SharedReg683_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg683_out;
SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg633_out;
SharedReg635_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg635_out;
SharedReg649_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg649_out;
SharedReg740_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg740_out;
SharedReg748_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg748_out;
SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg654_out;
SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg651_out;
SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg673_out;
SharedReg610_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg610_out;
SharedReg728_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg728_out;
SharedReg653_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg653_out;
SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg673_out;
   MUX_Product_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_36_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg674_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg685_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg671_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg719_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg665_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg737_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg614_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg681_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg677_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg646_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg720_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg611_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg666_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg683_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg633_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg635_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg649_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg740_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg748_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg636_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg610_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg728_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg653_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg673_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_4 => SharedReg658_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg654_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg716_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg657_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg691_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg651_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_2_impl_1_LUT_out,
                 oMux => MUX_Product_2_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product_3_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product_3_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_3_impl_out,
                 X => Delay1No4_out_to_Product_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product_3_impl_parent_implementedSystem_port_1_cast);

SharedReg423_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg423_out;
SharedReg341_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg345_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg351_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg351_out;
SharedReg349_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg349_out;
SharedReg356_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg356_out;
SharedReg357_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg357_out;
Delay91No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_8_cast <= Delay91No1_out;
SharedReg359_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg359_out;
SharedReg363_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg363_out;
SharedReg364_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg364_out;
SharedReg370_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg370_out;
SharedReg367_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg367_out;
SharedReg375_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg375_out;
SharedReg376_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg376_out;
SharedReg381_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg381_out;
SharedReg380_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg380_out;
SharedReg385_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg385_out;
SharedReg391_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg391_out;
SharedReg392_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg392_out;
SharedReg394_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg394_out;
SharedReg398_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg398_out;
SharedReg397_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg397_out;
SharedReg399_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg399_out;
SharedReg403_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg403_out;
SharedReg405_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg405_out;
SharedReg412_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg412_out;
SharedReg413_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg413_out;
SharedReg414_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg414_out;
SharedReg425_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg425_out;
SharedReg430_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg430_out;
SharedReg427_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg427_out;
SharedReg432_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg432_out;
SharedReg436_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg436_out;
Delay211No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_35_cast <= Delay211No1_out;
SharedReg442_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg442_out;
SharedReg448_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg448_out;
SharedReg447_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg447_out;
Delay67No2_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_39_cast <= Delay67No2_out;
SharedReg453_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg453_out;
SharedReg452_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg452_out;
SharedReg456_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg456_out;
Delay38No_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_43_cast <= Delay38No_out;
SharedReg460_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg460_out;
Delay75No3_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_45_cast <= Delay75No3_out;
SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg464_out;
SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg464_out;
SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg473_out;
SharedReg474_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg474_out;
SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg473_out;
   MUX_Product_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_50_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg423_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg364_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg370_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg367_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg375_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg376_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg381_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg380_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg385_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg391_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg392_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg345_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg394_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg398_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg397_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg399_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg403_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg405_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg412_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg413_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg414_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg425_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg351_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg430_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg427_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg432_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg436_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay211No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg442_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg448_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg447_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => Delay67No2_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg453_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg349_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg452_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg456_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => Delay38No_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg460_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay75No3_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg464_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg474_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg473_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg356_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg357_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay91No1_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg359_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg363_out_to_MUX_Product_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_3_impl_0_LUT_out,
                 oMux => MUX_Product_3_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_3_impl_0_out,
                 Y => Delay1No4_out);

SharedReg633_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg633_out;
SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg697_out;
SharedReg622_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg622_out;
SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg632_out;
SharedReg710_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg710_out;
SharedReg735_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg735_out;
SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg653_out;
SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg707_out;
SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg653_out;
SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg653_out;
SharedReg676_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg676_out;
SharedReg655_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg655_out;
SharedReg648_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg648_out;
SharedReg646_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg646_out;
SharedReg715_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg715_out;
SharedReg614_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg614_out;
SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg706_out;
SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg632_out;
SharedReg647_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg647_out;
SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg642_out;
SharedReg687_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg687_out;
SharedReg672_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg672_out;
SharedReg695_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg695_out;
SharedReg656_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg656_out;
SharedReg680_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg680_out;
SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg707_out;
SharedReg637_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg637_out;
SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg642_out;
SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg706_out;
SharedReg725_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg725_out;
SharedReg700_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg700_out;
SharedReg636_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg636_out;
SharedReg729_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg729_out;
SharedReg739_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg739_out;
Delay225No_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_35_cast <= Delay225No_out;
Delay135No3_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_36_cast <= Delay135No3_out;
SharedReg664_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg664_out;
SharedReg704_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg704_out;
SharedReg724_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg724_out;
SharedReg679_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg679_out;
SharedReg698_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg698_out;
SharedReg743_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg743_out;
SharedReg701_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg701_out;
SharedReg721_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg721_out;
SharedReg692_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg692_out;
SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg653_out;
SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg697_out;
SharedReg612_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg612_out;
SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg653_out;
SharedReg730_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg730_out;
   MUX_Product_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_50_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg633_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg676_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg655_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg648_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg646_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg715_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg614_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg647_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg622_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg687_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg672_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg695_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg656_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg680_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg637_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg642_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg706_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg725_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg632_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg700_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg636_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg729_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg739_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay225No_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => Delay135No3_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg664_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg704_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg724_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg679_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg710_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg698_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg743_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg701_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg721_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg692_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg697_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg612_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg730_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg735_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg707_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg653_out_to_MUX_Product_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_3_impl_1_LUT_out,
                 oMux => MUX_Product_3_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_3_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product1_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product1_2_impl_out,
                 X => Delay1No6_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast);

Delay13No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast <= Delay13No_out;
SharedReg344_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg342_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg374_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg374_out;
Delay88No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast <= Delay88No1_out;
Delay90No2_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast <= Delay90No2_out;
SharedReg389_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg389_out;
SharedReg401_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg401_out;
SharedReg402_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg402_out;
SharedReg408_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg408_out;
Delay169No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast <= Delay169No_out;
SharedReg411_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg411_out;
Delay61No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast <= Delay61No_out;
SharedReg416_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg416_out;
SharedReg417_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg417_out;
SharedReg421_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg421_out;
SharedReg422_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg422_out;
SharedReg429_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg429_out;
SharedReg433_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg433_out;
Delay17No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_20_cast <= Delay17No1_out;
SharedReg438_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg438_out;
SharedReg443_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg443_out;
SharedReg441_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg441_out;
SharedReg457_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg457_out;
SharedReg469_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg469_out;
SharedReg472_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg472_out;
   MUX_Product1_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay13No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay169No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg411_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay61No_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg416_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg417_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg421_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg422_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg429_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg433_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay17No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg438_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg443_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg441_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg457_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg469_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg472_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg374_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay88No1_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay90No2_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg389_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg401_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg402_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg408_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product1_2_impl_0_LUT_out,
                 oMux => MUX_Product1_2_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1_2_impl_0_out,
                 Y => Delay1No6_out);

SharedReg675_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg675_out;
SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg655_out;
SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg655_out;
SharedReg632_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg632_out;
SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg673_out;
SharedReg628_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg628_out;
SharedReg745_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg745_out;
SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg676_out;
SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg676_out;
SharedReg677_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg677_out;
SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg653_out;
Delay122No1_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast <= Delay122No1_out;
SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg654_out;
SharedReg683_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg683_out;
SharedReg728_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg728_out;
SharedReg688_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg688_out;
SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg654_out;
SharedReg742_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg742_out;
SharedReg697_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg697_out;
SharedReg696_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg696_out;
SharedReg684_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg684_out;
SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg673_out;
SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg653_out;
SharedReg698_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg698_out;
SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg653_out;
SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg673_out;
   MUX_Product1_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_26_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg675_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay122No1_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg683_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg728_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg688_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg654_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg742_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg697_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg696_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg655_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg684_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg698_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg653_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_3 => SharedReg632_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg673_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg628_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg745_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg676_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg677_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product1_2_impl_1_LUT_out,
                 oMux => MUX_Product1_2_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1_2_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product11_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_4_impl_out,
                 X => Delay1No8_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg355_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg355_out;
SharedReg361_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg361_out;
SharedReg378_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg378_out;
SharedReg407_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg428_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg428_out;
SharedReg435_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg435_out;
SharedReg450_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg450_out;
SharedReg454_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg454_out;
SharedReg458_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg458_out;
SharedReg465_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg465_out;
SharedReg468_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg468_out;
   MUX_Product11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg355_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg361_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg468_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg378_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg428_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg435_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg450_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg454_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg458_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg465_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product11_4_impl_0_LUT_out,
                 oMux => MUX_Product11_4_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_0_out,
                 Y => Delay1No8_out);

SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg659_out;
SharedReg682_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg682_out;
SharedReg689_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg689_out;
SharedReg727_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg727_out;
SharedReg733_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg733_out;
SharedReg663_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg663_out;
SharedReg660_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg660_out;
SharedReg654_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg654_out;
SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg659_out;
SharedReg741_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg741_out;
SharedReg673_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg673_out;
   MUX_Product11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg682_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg673_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg689_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg727_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg733_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg663_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg660_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg654_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg659_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg741_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product11_4_impl_1_LUT_out,
                 oMux => MUX_Product11_4_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No10_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => Delay1No10_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Sum10_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_0_impl_out,
                 X => Delay1No12_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg66_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg84_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg621_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg621_out;
SharedReg1_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg285_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg57_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg57_out;
SharedReg619_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg619_out;
SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg614_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg632_out;
SharedReg115_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg115_out;
SharedReg633_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg633_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg608_out;
SharedReg173_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg173_out;
SharedReg60_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg60_out;
SharedReg246_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg246_out;
SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg610_out;
SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg174_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg632_out;
SharedReg478_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg478_out;
SharedReg128_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg614_out;
SharedReg305_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg305_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg608_out;
SharedReg234_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg234_out;
SharedReg242_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg242_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg608_out;
SharedReg662_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg662_out;
SharedReg301_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg301_out;
SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg8_out;
SharedReg192_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg192_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg608_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg632_out;
SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg697_out;
SharedReg14_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg14_out;
SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg610_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg608_out;
SharedReg15_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg15_out;
SharedReg74_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg74_out;
SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg23_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg632_out;
SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg653_out;
SharedReg710_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg710_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg632_out;
SharedReg187_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg187_out;
SharedReg296_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg296_out;
SharedReg188_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg188_out;
SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg697_out;
SharedReg254_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg254_out;
SharedReg130_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg130_out;
SharedReg199_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg199_out;
SharedReg674_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg674_out;
SharedReg26_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg26_out;
SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg632_out;
SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg653_out;
SharedReg722_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg722_out;
SharedReg709_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg709_out;
SharedReg89_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg89_out;
SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg608_out;
   MUX_Sum10_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg115_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg633_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg173_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg60_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg246_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg478_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg84_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg305_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg234_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg242_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg662_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg301_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg621_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg192_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg14_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg610_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg15_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg74_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg710_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg187_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg296_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg188_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg697_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg254_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg130_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg285_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg199_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg674_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg26_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg653_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg722_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg709_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg89_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg608_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg57_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg619_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg614_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg632_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_0_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_0_impl_0_out,
                 Y => Delay1No12_out);

SharedReg329_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg45_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg45_out;
SharedReg28_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg499_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg499_out;
Delay590No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast <= Delay590No_out;
SharedReg279_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg279_out;
Delay591No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast <= Delay591No_out;
SharedReg509_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg509_out;
SharedReg503_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg503_out;
SharedReg485_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg485_out;
Delay597No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast <= Delay597No_out;
SharedReg515_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg515_out;
SharedReg512_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg512_out;
Delay603No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast <= Delay603No_out;
SharedReg55_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg55_out;
SharedReg208_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg208_out;
SharedReg513_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg513_out;
Delay546No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast <= Delay546No_out;
SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg478_out;
SharedReg481_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg481_out;
SharedReg209_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg209_out;
SharedReg486_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg486_out;
SharedReg30_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg30_out;
SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg478_out;
SharedReg222_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg222_out;
SharedReg214_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg214_out;
SharedReg493_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg493_out;
SharedReg574_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg574_out;
SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg152_out;
SharedReg111_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg111_out;
SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg264_out;
SharedReg482_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg482_out;
SharedReg487_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg487_out;
SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg479_out;
SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg105_out;
SharedReg517_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg517_out;
SharedReg553_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg553_out;
SharedReg326_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg326_out;
SharedReg39_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg39_out;
SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg93_out;
SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg518_out;
SharedReg558_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg558_out;
SharedReg504_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg504_out;
SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg479_out;
SharedReg155_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg155_out;
SharedReg161_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg161_out;
SharedReg272_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg272_out;
SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg518_out;
SharedReg205_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg205_out;
SharedReg327_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg327_out;
SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg261_out;
SharedReg502_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg502_out;
SharedReg315_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg315_out;
SharedReg480_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg480_out;
SharedReg508_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg508_out;
SharedReg497_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg497_out;
SharedReg557_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg557_out;
SharedReg44_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg44_out;
SharedReg491_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg491_out;
   MUX_Sum10_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg45_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay597No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg515_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg512_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay603No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg55_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg208_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg513_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay546No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg481_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg28_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg209_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg486_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg30_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg478_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg222_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg214_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg493_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg574_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg111_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg499_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg482_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg487_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg517_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg553_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg326_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg39_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => Delay590No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg558_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg504_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg479_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg155_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg161_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg272_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg518_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg205_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg327_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg279_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg502_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg315_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg480_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg508_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg497_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg557_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg44_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg491_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => Delay591No_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg509_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg503_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg485_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_0_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_0_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Sum10_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_1_impl_out,
                 X => Delay1No14_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast);

SharedReg138_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg138_out;
SharedReg228_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg228_out;
Delay134No1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast <= Delay134No1_out;
SharedReg_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg_out;
SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg608_out;
SharedReg670_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg670_out;
SharedReg655_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg655_out;
SharedReg694_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg694_out;
SharedReg12_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg12_out;
SharedReg245_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg245_out;
SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg673_out;
SharedReg240_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg240_out;
SharedReg660_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg660_out;
SharedReg478_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg478_out;
SharedReg639_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg639_out;
SharedReg229_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg229_out;
SharedReg230_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg230_out;
SharedReg78_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg78_out;
SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg175_out;
SharedReg4_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg4_out;
SharedReg638_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg638_out;
SharedReg133_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg133_out;
SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg673_out;
SharedReg251_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg251_out;
SharedReg637_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg637_out;
SharedReg191_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg191_out;
SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg697_out;
SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg632_out;
SharedReg129_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg129_out;
SharedReg714_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg714_out;
SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg9_out;
SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg673_out;
SharedReg661_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg661_out;
SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg699_out;
SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg632_out;
SharedReg705_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg705_out;
SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg697_out;
SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg608_out;
SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg75_out;
SharedReg69_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg69_out;
SharedReg728_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg728_out;
SharedReg678_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg678_out;
SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg699_out;
SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg79_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg296_out;
SharedReg253_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg253_out;
SharedReg653_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg653_out;
SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg608_out;
SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg136_out;
SharedReg237_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg237_out;
SharedReg77_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg77_out;
SharedReg636_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg636_out;
SharedReg298_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg298_out;
SharedReg195_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg195_out;
SharedReg131_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg131_out;
SharedReg299_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg299_out;
SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg673_out;
SharedReg82_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg82_out;
   MUX_Sum10_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg138_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg240_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg660_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg478_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg639_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg229_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg230_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg78_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg4_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => Delay134No1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg638_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg133_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg251_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg637_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg191_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg129_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg714_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg661_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg632_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg705_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg697_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg69_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg728_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg678_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg699_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg253_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg653_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg608_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg670_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg237_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg77_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg636_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg298_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg195_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg131_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg299_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg673_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg82_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg655_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg694_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg12_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg245_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_1_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_1_impl_0_out,
                 Y => Delay1No14_out);

SharedReg83_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg335_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg335_out;
SharedReg488_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg488_out;
SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg225_out;
SharedReg494_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg494_out;
SharedReg487_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg487_out;
SharedReg579_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg579_out;
Delay249No1_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast <= Delay249No1_out;
SharedReg97_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg97_out;
SharedReg90_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg90_out;
SharedReg519_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg519_out;
SharedReg207_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg207_out;
SharedReg505_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg505_out;
SharedReg543_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg543_out;
SharedReg501_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg501_out;
SharedReg110_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg110_out;
SharedReg220_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg220_out;
SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg257_out;
SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg165_out;
SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg221_out;
SharedReg596_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg596_out;
SharedReg311_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg311_out;
SharedReg546_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg546_out;
SharedReg490_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg490_out;
SharedReg312_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg312_out;
SharedReg492_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg492_out;
SharedReg259_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg259_out;
SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg478_out;
SharedReg585_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg585_out;
SharedReg318_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg318_out;
SharedReg521_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg521_out;
SharedReg223_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg223_out;
SharedReg565_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg565_out;
Delay358No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast <= Delay358No_out;
Delay339No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast <= Delay339No_out;
SharedReg549_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg549_out;
SharedReg516_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg516_out;
SharedReg550_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg550_out;
SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg478_out;
SharedReg153_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg153_out;
SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg40_out;
SharedReg527_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg527_out;
SharedReg536_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg536_out;
SharedReg566_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg566_out;
SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg32_out;
SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg271_out;
SharedReg87_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg87_out;
SharedReg583_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg583_out;
SharedReg486_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg486_out;
SharedReg320_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg320_out;
SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg106_out;
SharedReg148_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg148_out;
SharedReg578_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg578_out;
SharedReg42_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg42_out;
SharedReg37_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg37_out;
SharedReg100_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg100_out;
SharedReg266_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg266_out;
SharedReg485_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg485_out;
SharedReg149_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg149_out;
   MUX_Sum10_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg519_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg207_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg505_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg543_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg501_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg110_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg220_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg488_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg596_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg311_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg546_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg490_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg312_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg492_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg259_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg585_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg318_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg521_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg223_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg565_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay358No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay339No_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg549_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg516_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg550_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg478_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg153_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg494_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg527_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg536_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg566_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg87_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg583_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg486_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg320_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg487_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg148_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg578_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg42_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg37_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg100_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg266_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg485_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg149_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg579_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay249No1_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg97_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg90_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_1_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_1_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Sum10_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_2_impl_out,
                 X => Delay1No16_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast);

SharedReg699_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg283_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg283_out;
SharedReg282_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg282_out;
SharedReg701_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg701_out;
SharedReg169_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg169_out;
SharedReg56_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg56_out;
SharedReg727_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg727_out;
SharedReg190_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg190_out;
SharedReg171_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg171_out;
SharedReg668_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg668_out;
SharedReg115_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg115_out;
SharedReg675_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg675_out;
SharedReg58_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg58_out;
SharedReg720_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg720_out;
SharedReg634_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg634_out;
SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg124_out;
SharedReg658_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg658_out;
SharedReg287_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg287_out;
SharedReg3_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg3_out;
SharedReg288_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg288_out;
SharedReg669_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg669_out;
SharedReg5_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg5_out;
SharedReg656_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg656_out;
SharedReg662_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg662_out;
SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg186_out;
SharedReg231_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg231_out;
SharedReg63_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg63_out;
SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg632_out;
SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg635_out;
SharedReg119_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg119_out;
SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg632_out;
SharedReg697_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg697_out;
SharedReg293_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg293_out;
SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg10_out;
SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg193_out;
SharedReg661_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg661_out;
SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg635_out;
SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg632_out;
SharedReg121_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg121_out;
SharedReg183_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg183_out;
SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg673_out;
SharedReg729_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg729_out;
SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg632_out;
SharedReg64_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg64_out;
SharedReg236_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg236_out;
SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg18_out;
SharedReg71_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg71_out;
SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg673_out;
SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg632_out;
SharedReg702_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg702_out;
SharedReg76_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg76_out;
SharedReg730_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg730_out;
SharedReg256_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg256_out;
SharedReg137_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg137_out;
SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg20_out;
SharedReg21_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg27_out;
SharedReg238_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg238_out;
SharedReg633_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg633_out;
   MUX_Sum10_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg283_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg115_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg675_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg58_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg720_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg634_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg658_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg287_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg3_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg288_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg282_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg669_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg5_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg656_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg662_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg231_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg63_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg119_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg701_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg697_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg293_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg661_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg635_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg121_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg183_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg169_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg729_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg64_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg236_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg71_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg673_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg632_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg702_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg56_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg76_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg730_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg256_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg137_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg21_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg27_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg238_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg633_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg727_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg190_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg171_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg668_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_2_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_2_impl_0_out,
                 Y => Delay1No16_out);

SharedReg524_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg524_out;
SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg51_out;
SharedReg52_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg539_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg539_out;
SharedReg53_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg53_out;
SharedReg54_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg54_out;
SharedReg538_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg538_out;
SharedReg29_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg29_out;
SharedReg280_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg280_out;
SharedReg542_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg542_out;
SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg219_out;
SharedReg573_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg573_out;
SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg163_out;
SharedReg510_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg510_out;
SharedReg599_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg599_out;
SharedReg323_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg323_out;
SharedReg535_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg535_out;
SharedReg164_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg164_out;
Delay607No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast <= Delay607No_out;
SharedReg276_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg276_out;
SharedReg517_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg517_out;
SharedReg331_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg331_out;
SharedReg598_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg598_out;
SharedReg576_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg576_out;
SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg263_out;
SharedReg332_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg332_out;
SharedReg160_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg160_out;
SharedReg522_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg522_out;
SharedReg580_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg580_out;
SharedReg102_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg102_out;
SharedReg553_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg553_out;
SharedReg572_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg572_out;
SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg269_out;
SharedReg104_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg104_out;
SharedReg145_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg145_out;
SharedReg607_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg607_out;
SharedReg526_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg526_out;
SharedReg532_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg532_out;
SharedReg333_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg333_out;
SharedReg49_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg49_out;
SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg547_out;
SharedReg594_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg594_out;
SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg547_out;
SharedReg50_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg50_out;
SharedReg98_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg98_out;
SharedReg212_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg212_out;
SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg265_out;
SharedReg511_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg511_out;
SharedReg577_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg577_out;
SharedReg507_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg507_out;
SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg261_out;
SharedReg588_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg588_out;
SharedReg200_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg200_out;
SharedReg206_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg206_out;
SharedReg95_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg95_out;
SharedReg322_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg322_out;
SharedReg201_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg201_out;
SharedReg328_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg328_out;
SharedReg541_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg541_out;
   MUX_Sum10_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg524_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg573_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg510_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg599_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg323_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg535_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg164_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => Delay607No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg276_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg52_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg517_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg331_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg598_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg576_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg332_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg160_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg522_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg580_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg102_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg539_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg553_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg572_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg104_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg145_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg607_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg526_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg532_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg333_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg49_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg53_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg594_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg547_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg50_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg98_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg212_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg511_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg577_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg507_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg54_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg588_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg200_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg206_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg95_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg322_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg201_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg328_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg541_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg538_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg29_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg280_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg542_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_2_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_2_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Sum10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_3_impl_out,
                 X => Delay1No18_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg244_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg178_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg178_out;
SharedReg226_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg72_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg72_out;
SharedReg675_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg675_out;
SharedReg674_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg674_out;
SharedReg123_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg170_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg170_out;
SharedReg114_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg114_out;
SharedReg2_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg2_out;
SharedReg239_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg239_out;
SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg518_out;
SharedReg286_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg286_out;
SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg518_out;
SharedReg132_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg132_out;
SharedReg73_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg73_out;
SharedReg184_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg184_out;
SharedReg543_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg543_out;
SharedReg633_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg633_out;
SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg185_out;
SharedReg295_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg295_out;
SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg727_out;
SharedReg659_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg659_out;
SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg727_out;
SharedReg176_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg176_out;
SharedReg300_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg300_out;
SharedReg243_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg243_out;
SharedReg734_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg734_out;
SharedReg306_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg306_out;
SharedReg13_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg13_out;
SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg181_out;
SharedReg709_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg709_out;
SharedReg232_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg232_out;
SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg727_out;
SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg177_out;
SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg653_out;
SharedReg235_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg235_out;
SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg135_out;
SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg673_out;
SharedReg68_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg68_out;
SharedReg666_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg666_out;
SharedReg248_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg248_out;
SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg653_out;
SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg673_out;
SharedReg127_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg127_out;
SharedReg608_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg608_out;
SharedReg16_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg16_out;
SharedReg249_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg249_out;
SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg11_out;
SharedReg130_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg130_out;
SharedReg80_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg80_out;
SharedReg297_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg297_out;
SharedReg632_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg632_out;
SharedReg654_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg654_out;
SharedReg310_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg310_out;
SharedReg616_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg616_out;
SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg653_out;
SharedReg744_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg744_out;
SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg727_out;
   MUX_Sum10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg178_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg239_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg286_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg518_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg132_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg73_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg184_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg543_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg633_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg226_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg295_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg659_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg176_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg300_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg243_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg734_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg306_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg13_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg72_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg709_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg232_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg235_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg68_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg675_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg666_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg248_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg673_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg127_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg608_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg16_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg249_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg130_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg674_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg80_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg297_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg632_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg654_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg310_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg616_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg653_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg744_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg727_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg123_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg170_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg114_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg2_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_3_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_3_impl_0_out,
                 Y => Delay1No18_out);

SharedReg202_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg267_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg267_out;
SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg107_out;
SharedReg262_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg568_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg601_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg601_out;
SharedReg96_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg96_out;
SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg337_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg337_out;
SharedReg109_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg109_out;
SharedReg91_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg91_out;
SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg583_out;
SharedReg47_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg47_out;
SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg583_out;
SharedReg196_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg196_out;
SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg33_out;
SharedReg144_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg144_out;
SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg518_out;
SharedReg555_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg555_out;
SharedReg34_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg34_out;
SharedReg151_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg151_out;
SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg583_out;
SharedReg584_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg584_out;
SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg583_out;
SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg159_out;
SharedReg258_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg258_out;
SharedReg317_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg317_out;
SharedReg592_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg592_out;
SharedReg252_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg252_out;
SharedReg210_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg210_out;
SharedReg38_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg38_out;
SharedReg567_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg567_out;
SharedReg103_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg103_out;
SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg518_out;
SharedReg48_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg48_out;
SharedReg531_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg531_out;
SharedReg215_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg215_out;
SharedReg85_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg85_out;
SharedReg544_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg544_out;
SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg270_out;
SharedReg578_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg578_out;
SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg86_out;
SharedReg484_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg484_out;
SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg518_out;
SharedReg211_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg211_out;
SharedReg562_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg562_out;
SharedReg319_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg319_out;
SharedReg314_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg314_out;
SharedReg334_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg334_out;
SharedReg94_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg94_out;
SharedReg255_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg255_out;
SharedReg36_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg36_out;
SharedReg543_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg543_out;
SharedReg591_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg591_out;
SharedReg142_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg142_out;
SharedReg509_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg509_out;
Delay103No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast <= Delay103No_out;
SharedReg540_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg540_out;
SharedReg554_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg554_out;
   MUX_Sum10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg267_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg91_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg47_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg196_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg144_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg555_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg34_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg151_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg584_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg583_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg258_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg317_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg592_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg252_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg210_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg262_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg38_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg567_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg103_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg48_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg531_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg215_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg85_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg544_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg568_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg578_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg484_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg518_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg211_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg562_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg319_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg314_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg334_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg94_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg601_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg255_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg36_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg543_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg591_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg142_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg509_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => Delay103No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg540_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg554_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg96_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg337_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg109_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_3_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_3_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Sum11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Sum11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Sum11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum11_0_impl_out,
                 X => Delay1No20_out_to_Sum11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Sum11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg22_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg228_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg228_out;
SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg608_out;
SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg610_out;
SharedReg284_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg699_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg699_out;
SharedReg618_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg618_out;
SharedReg179_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg179_out;
SharedReg679_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg679_out;
SharedReg116_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg116_out;
SharedReg6_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg290_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg290_out;
SharedReg58_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg58_out;
SharedReg117_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg117_out;
SharedReg291_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg291_out;
SharedReg67_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg67_out;
SharedReg241_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg241_out;
SharedReg233_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg233_out;
SharedReg704_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg704_out;
SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg610_out;
SharedReg197_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg197_out;
SharedReg61_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg61_out;
SharedReg518_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg518_out;
SharedReg125_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg125_out;
SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg610_out;
SharedReg292_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg292_out;
SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg616_out;
SharedReg715_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg715_out;
SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg608_out;
SharedReg247_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg247_out;
SharedReg120_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg120_out;
SharedReg198_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg198_out;
SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg653_out;
SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg616_out;
SharedReg625_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg625_out;
SharedReg134_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg134_out;
SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg653_out;
SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg608_out;
SharedReg182_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg182_out;
SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg697_out;
SharedReg126_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg126_out;
SharedReg70_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg70_out;
SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg697_out;
SharedReg307_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg307_out;
SharedReg303_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg303_out;
SharedReg141_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg141_out;
SharedReg304_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg304_out;
SharedReg717_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg717_out;
SharedReg308_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg308_out;
SharedReg19_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg19_out;
SharedReg250_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg250_out;
SharedReg25_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg25_out;
SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg697_out;
SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg653_out;
SharedReg189_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg189_out;
SharedReg65_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg65_out;
SharedReg643_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg643_out;
SharedReg609_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg609_out;
SharedReg17_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg17_out;
   MUX_Sum11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg290_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg58_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg117_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg291_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg67_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg241_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg233_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg704_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg197_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg61_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg518_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg125_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg292_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg715_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg247_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg610_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg120_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg198_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg616_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg625_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg134_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg608_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg182_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg284_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg126_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg70_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg307_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg303_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg141_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg304_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg717_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg308_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg19_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg699_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg250_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg25_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg697_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg653_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg189_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg65_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg643_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg609_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg17_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg618_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg179_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg679_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg116_out_to_MUX_Sum11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum11_0_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum11_0_impl_0_out,
                 Y => Delay1No20_out);

SharedReg202_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg224_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg224_out;
SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg551_out;
SharedReg570_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg168_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg168_out;
SharedReg491_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg491_out;
SharedReg484_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg484_out;
SharedReg157_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg157_out;
SharedReg537_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg537_out;
SharedReg218_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg218_out;
SharedReg213_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg213_out;
SharedReg46_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg281_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg281_out;
SharedReg338_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg338_out;
SharedReg274_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg274_out;
SharedReg158_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg158_out;
SharedReg324_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg324_out;
SharedReg330_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg330_out;
SharedReg569_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg569_out;
SharedReg582_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg582_out;
SharedReg139_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg139_out;
SharedReg277_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg277_out;
SharedReg583_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg583_out;
SharedReg101_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg101_out;
SharedReg514_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg514_out;
SharedReg166_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg166_out;
SharedReg504_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg504_out;
SharedReg498_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg498_out;
SharedReg545_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg545_out;
SharedReg102_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg102_out;
SharedReg112_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg112_out;
SharedReg31_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg31_out;
SharedReg600_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg600_out;
SharedReg552_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg552_out;
SharedReg500_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg500_out;
SharedReg92_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg92_out;
SharedReg575_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg575_out;
SharedReg483_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg483_out;
SharedReg278_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg278_out;
SharedReg506_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg506_out;
SharedReg216_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg216_out;
SharedReg154_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg154_out;
SharedReg523_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg523_out;
SharedReg260_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg260_out;
SharedReg35_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg35_out;
SharedReg313_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg313_out;
SharedReg265_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg265_out;
SharedReg495_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg495_out;
SharedReg147_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg147_out;
SharedReg99_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg99_out;
SharedReg321_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg321_out;
SharedReg88_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg88_out;
SharedReg528_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg528_out;
SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg551_out;
SharedReg43_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg43_out;
SharedReg167_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg167_out;
SharedReg566_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg566_out;
SharedReg560_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg560_out;
SharedReg217_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg217_out;
   MUX_Sum11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg224_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg213_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg281_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg338_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg274_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg158_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg324_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg330_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg569_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg582_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg139_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg277_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg583_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg101_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg514_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg166_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg504_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg498_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg545_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg102_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg570_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg112_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg31_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg600_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg552_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg500_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg92_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg575_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg483_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg278_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg506_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg168_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg216_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg154_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg523_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg260_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg35_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg313_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg265_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg495_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg147_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg99_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg491_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg321_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg88_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg528_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg551_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg43_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg167_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg566_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg560_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg217_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg484_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg157_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg537_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg218_out_to_MUX_Sum11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum11_0_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum11_0_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Sum11_5_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Sum11_5_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Sum11_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum11_5_impl_out,
                 X => Delay1No22_out_to_Sum11_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Sum11_5_impl_parent_implementedSystem_port_1_cast);

SharedReg289_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg289_out;
SharedReg675_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg675_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg727_out;
SharedReg227_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg227_out;
SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg728_out;
SharedReg113_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg113_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg727_out;
SharedReg667_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg667_out;
SharedReg172_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg172_out;
SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg728_out;
SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg738_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg727_out;
SharedReg637_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg637_out;
SharedReg747_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg747_out;
SharedReg59_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg59_out;
SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg673_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg727_out;
SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg673_out;
SharedReg180_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg180_out;
SharedReg128_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg128_out;
SharedReg732_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg732_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg727_out;
SharedReg62_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg62_out;
SharedReg7_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg7_out;
SharedReg118_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg118_out;
SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg673_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg727_out;
SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg673_out;
SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg738_out;
SharedReg746_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg746_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg727_out;
SharedReg735_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg735_out;
SharedReg679_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg679_out;
SharedReg645_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg645_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg727_out;
SharedReg731_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg731_out;
SharedReg302_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg302_out;
SharedReg194_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg194_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg727_out;
SharedReg303_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg303_out;
SharedReg18_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg18_out;
SharedReg742_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg742_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg727_out;
SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg673_out;
SharedReg294_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg294_out;
SharedReg24_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg24_out;
SharedReg736_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg736_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg727_out;
SharedReg20_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg20_out;
SharedReg81_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg81_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg727_out;
SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg727_out;
SharedReg640_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg640_out;
   MUX_Sum11_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg289_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg675_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg637_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg747_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg59_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg180_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg128_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg732_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg62_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg7_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg118_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg738_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg227_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg746_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg735_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg679_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg645_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg731_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg302_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg194_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg303_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg18_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg742_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg673_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg294_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg728_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg24_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg736_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg20_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg81_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg640_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg113_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg727_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg667_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg172_out_to_MUX_Sum11_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum11_5_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum11_5_impl_0_out,
                 Y => Delay1No22_out);

SharedReg156_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg156_out;
SharedReg571_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg571_out;
SharedReg561_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg561_out;
SharedReg336_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg336_out;
SharedReg605_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg605_out;
SharedReg589_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg589_out;
SharedReg108_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg108_out;
SharedReg602_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg602_out;
SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg564_out;
SharedReg273_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg273_out;
SharedReg606_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg606_out;
SharedReg594_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg594_out;
SharedReg563_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg563_out;
Delay296No_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_14_cast <= Delay296No_out;
SharedReg595_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg595_out;
SharedReg275_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg275_out;
SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg518_out;
SharedReg587_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg587_out;
SharedReg543_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg543_out;
SharedReg150_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg150_out;
SharedReg203_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg203_out;
SharedReg581_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg581_out;
SharedReg530_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg530_out;
SharedReg268_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg268_out;
SharedReg325_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg325_out;
SharedReg214_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg214_out;
SharedReg478_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg478_out;
SharedReg525_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg525_out;
SharedReg583_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg583_out;
SharedReg489_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg489_out;
SharedReg586_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg586_out;
SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg518_out;
SharedReg496_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg496_out;
Delay351No2_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_34_cast <= Delay351No2_out;
SharedReg596_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg596_out;
SharedReg559_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg559_out;
SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg600_out;
SharedReg590_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg590_out;
SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg564_out;
SharedReg146_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg146_out;
SharedReg140_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg140_out;
SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg600_out;
SharedReg603_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg603_out;
SharedReg533_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg533_out;
SharedReg32_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg32_out;
SharedReg204_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg204_out;
SharedReg597_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg597_out;
SharedReg534_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg534_out;
SharedReg548_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg548_out;
SharedReg41_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg41_out;
SharedReg309_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg309_out;
SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg529_out;
SharedReg593_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg593_out;
SharedReg520_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg520_out;
SharedReg316_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg316_out;
SharedReg143_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg143_out;
SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg529_out;
SharedReg604_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg604_out;
SharedReg556_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg556_out;
   MUX_Sum11_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg156_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg571_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg606_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg594_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg563_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay296No_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg595_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg275_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg587_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg543_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg150_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg561_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg203_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg581_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg530_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg268_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg325_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg214_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg478_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg525_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg583_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg489_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg336_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg586_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg518_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg496_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay351No2_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg596_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg559_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg590_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg146_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg605_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg140_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg600_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg603_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg533_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg32_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg204_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg597_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg534_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg548_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg41_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg589_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg309_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg593_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg520_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg316_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg143_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg529_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg604_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg556_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg108_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg602_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg564_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg273_out_to_MUX_Sum11_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum11_5_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum11_5_impl_1_out,
                 Y => Delay1No23_out);
   Y_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_0_IEEE,
                 X => Delay1No24_out);
Y_0 <= Y_0_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => Delay1No24_out);
   Y_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_1_IEEE,
                 X => Delay1No25_out);
Y_1 <= Y_1_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => Delay1No25_out);
   Y_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_2_IEEE,
                 X => Delay1No26_out);
Y_2 <= Y_2_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => Delay1No26_out);
   Y_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_3_IEEE,
                 X => Delay1No27_out);
Y_3 <= Y_3_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => Delay1No27_out);
   Y_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_4_IEEE,
                 X => Delay1No28_out);
Y_4 <= Y_4_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => Delay1No28_out);
   Y_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_5_IEEE,
                 X => Delay1No29_out);
Y_5 <= Y_5_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => Delay1No29_out);

   Delay546No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => Delay546No_out);

   Delay590No_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => Delay590No_out);

   Delay591No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => Delay591No_out);

   Delay597No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => Delay597No_out);

   Delay603No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => Delay603No_out);

   Delay607No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => Delay607No_out);

   Delay18No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => Delay18No_out);

   Delay13No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => Delay13No_out);

   Delay102No_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => Delay102No_out);

   Delay77No1_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => Delay77No1_out);

   Delay91No1_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => Delay91No1_out);

   Delay101No_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => Delay101No_out);

   Delay107No_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay107No_out);

   Delay91No2_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => Delay91No2_out);

   Delay138No_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => Delay138No_out);

   Delay88No1_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => Delay88No1_out);

   Delay90No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => Delay90No2_out);

   Delay111No_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => Delay111No_out);

   Delay19No3_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => Delay19No3_out);

   Delay109No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => Delay109No_out);

   Delay169No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => Delay169No_out);

   Delay61No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => Delay61No_out);

   Delay65No1_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => Delay65No1_out);

   Delay322No1_instance: Delay_34_DelayLength_70_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=70 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => Delay322No1_out);

   Delay323No2_instance: Delay_34_DelayLength_160_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=160 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => Delay323No2_out);

   Delay161No_instance: Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=105 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => Delay161No_out);

   Delay17No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => Delay17No1_out);

   Delay211No1_instance: Delay_34_DelayLength_146_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=146 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => Delay211No1_out);

   Delay67No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => Delay67No2_out);

   Delay278No_instance: Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=103 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => Delay278No_out);

   Delay38No_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => Delay38No_out);

   Delay76No1_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => Delay76No1_out);

   Delay75No3_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => Delay75No3_out);

   Delay95No_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => Delay95No_out);

   Delay52No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => Delay52No2_out);

   Delay55No1_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => Delay55No1_out);

   Delay249No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => Delay249No1_out);

   Delay296No_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => Delay296No_out);

   Delay339No_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => Delay339No_out);

   Delay358No_instance: Delay_34_DelayLength_66_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=66 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => Delay358No_out);

   Delay351No2_instance: Delay_34_DelayLength_101_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=101 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => Delay351No2_out);

   Delay103No_instance: Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=103 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => Delay103No_out);

   Delay122No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => Delay122No1_out);

   Delay225No_instance: Delay_34_DelayLength_115_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=115 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => Delay225No_out);

   Delay135No3_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => Delay135No3_out);

   Delay266No1_instance: Delay_34_DelayLength_154_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=154 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => Delay266No1_out);

   Delay288No_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => Delay288No_out);

   Delay134No1_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => Delay134No1_out);

   MUX_Product_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_0_impl_0_LUT_out);

   MUX_Product_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_0_impl_1_LUT_out);

   MUX_Product_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_2_impl_0_LUT_out);

   MUX_Product_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_2_impl_1_LUT_out);

   MUX_Product_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_3_impl_0_LUT_out);

   MUX_Product_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_3_impl_1_LUT_out);

   MUX_Product1_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product1_2_impl_0_LUT_out);

   MUX_Product1_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product1_2_impl_1_LUT_out);

   MUX_Product11_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product11_4_impl_0_LUT_out);

   MUX_Product11_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product11_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_1_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_2_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_3_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_4_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_5_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant10_0_impl_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant12_0_impl_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant19_0_impl_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant20_0_impl_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant21_0_impl_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_88_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=88 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant22_0_impl_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant23_0_impl_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant24_0_impl_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_74_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=74 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant25_0_impl_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_86_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=86 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant29_0_impl_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant3_0_impl_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant32_0_impl_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant33_0_impl_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant34_0_impl_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_33_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=33 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_117_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=117 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_0_impl_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_2_impl_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_3_impl_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product1_2_impl_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_4_impl_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=59 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_141_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=141 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_0_impl_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_60_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=60 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_1_impl_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_2_impl_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_3_impl_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum11_0_impl_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_82_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=82 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum11_5_impl_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);
end architecture;

